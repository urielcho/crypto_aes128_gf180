* NGSPICE file created from user_project_wrapper.ext - technology: gf180mcuC

* Black-box entry subcircuit for aes128 abstract view
.subckt aes128 clk key[0] key[100] key[101] key[102] key[103] key[104] key[105] key[106]
+ key[107] key[108] key[109] key[10] key[110] key[111] key[112] key[113] key[114]
+ key[115] key[116] key[117] key[118] key[119] key[11] key[120] key[121] key[122]
+ key[123] key[124] key[125] key[126] key[127] key[12] key[13] key[14] key[15] key[16]
+ key[17] key[18] key[19] key[1] key[20] key[21] key[22] key[23] key[24] key[25] key[26]
+ key[27] key[28] key[29] key[2] key[30] key[31] key[32] key[33] key[34] key[35] key[36]
+ key[37] key[38] key[39] key[3] key[40] key[41] key[42] key[43] key[44] key[45] key[46]
+ key[47] key[48] key[49] key[4] key[50] key[51] key[52] key[53] key[54] key[55] key[56]
+ key[57] key[58] key[59] key[5] key[60] key[61] key[62] key[63] key[64] key[65] key[66]
+ key[67] key[68] key[69] key[6] key[70] key[71] key[72] key[73] key[74] key[75] key[76]
+ key[77] key[78] key[79] key[7] key[80] key[81] key[82] key[83] key[84] key[85] key[86]
+ key[87] key[88] key[89] key[8] key[90] key[91] key[92] key[93] key[94] key[95] key[96]
+ key[97] key[98] key[99] key[9] out[0] out[100] out[101] out[102] out[103] out[104]
+ out[105] out[106] out[107] out[108] out[109] out[10] out[110] out[111] out[112]
+ out[113] out[114] out[115] out[116] out[117] out[118] out[119] out[11] out[120]
+ out[121] out[122] out[123] out[124] out[125] out[126] out[127] out[12] out[13] out[14]
+ out[15] out[16] out[17] out[18] out[19] out[1] out[20] out[21] out[22] out[23] out[24]
+ out[25] out[26] out[27] out[28] out[29] out[2] out[30] out[31] out[32] out[33] out[34]
+ out[35] out[36] out[37] out[38] out[39] out[3] out[40] out[41] out[42] out[43] out[44]
+ out[45] out[46] out[47] out[48] out[49] out[4] out[50] out[51] out[52] out[53] out[54]
+ out[55] out[56] out[57] out[58] out[59] out[5] out[60] out[61] out[62] out[63] out[64]
+ out[65] out[66] out[67] out[68] out[69] out[6] out[70] out[71] out[72] out[73] out[74]
+ out[75] out[76] out[77] out[78] out[79] out[7] out[80] out[81] out[82] out[83] out[84]
+ out[85] out[86] out[87] out[88] out[89] out[8] out[90] out[91] out[92] out[93] out[94]
+ out[95] out[96] out[97] out[98] out[99] out[9] state[0] state[100] state[101] state[102]
+ state[103] state[104] state[105] state[106] state[107] state[108] state[109] state[10]
+ state[110] state[111] state[112] state[113] state[114] state[115] state[116] state[117]
+ state[118] state[119] state[11] state[120] state[121] state[122] state[123] state[124]
+ state[125] state[126] state[127] state[12] state[13] state[14] state[15] state[16]
+ state[17] state[18] state[19] state[1] state[20] state[21] state[22] state[23] state[24]
+ state[25] state[26] state[27] state[28] state[29] state[2] state[30] state[31] state[32]
+ state[33] state[34] state[35] state[36] state[37] state[38] state[39] state[3] state[40]
+ state[41] state[42] state[43] state[44] state[45] state[46] state[47] state[48]
+ state[49] state[4] state[50] state[51] state[52] state[53] state[54] state[55] state[56]
+ state[57] state[58] state[59] state[5] state[60] state[61] state[62] state[63] state[64]
+ state[65] state[66] state[67] state[68] state[69] state[6] state[70] state[71] state[72]
+ state[73] state[74] state[75] state[76] state[77] state[78] state[79] state[7] state[80]
+ state[81] state[82] state[83] state[84] state[85] state[86] state[87] state[88]
+ state[89] state[8] state[90] state[91] state[92] state[93] state[94] state[95] state[96]
+ state[97] state[98] state[99] state[9] vdd vss
.ends

.subckt user_project_wrapper io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10]
+ la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15]
+ la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20]
+ la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25]
+ la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30]
+ la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40]
+ la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50]
+ la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55]
+ la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60]
+ la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[6] la_oenb[7]
+ la_oenb[8] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2] vdd vss wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xaes128 wb_clk_i aes128/key[0] aes128/key[100] aes128/key[101] aes128/key[102] aes128/key[103]
+ aes128/key[104] aes128/key[105] aes128/key[106] aes128/key[107] aes128/key[108]
+ aes128/key[109] aes128/key[10] aes128/key[110] aes128/key[111] aes128/key[112] aes128/key[113]
+ aes128/key[114] aes128/key[115] aes128/key[116] aes128/key[117] aes128/key[118]
+ aes128/key[119] aes128/key[11] aes128/key[120] aes128/key[121] aes128/key[122] aes128/key[123]
+ aes128/key[124] aes128/key[125] aes128/key[126] aes128/key[127] aes128/key[12] aes128/key[13]
+ aes128/key[14] aes128/key[15] aes128/key[16] aes128/key[17] aes128/key[18] aes128/key[19]
+ aes128/key[1] aes128/key[20] aes128/key[21] aes128/key[22] aes128/key[23] aes128/key[24]
+ aes128/key[25] aes128/key[26] aes128/key[27] aes128/key[28] aes128/key[29] aes128/key[2]
+ aes128/key[30] aes128/key[31] aes128/key[32] aes128/key[33] aes128/key[34] aes128/key[35]
+ aes128/key[36] aes128/key[37] aes128/key[38] aes128/key[39] aes128/key[3] aes128/key[40]
+ aes128/key[41] aes128/key[42] aes128/key[43] aes128/key[44] aes128/key[45] aes128/key[46]
+ aes128/key[47] aes128/key[48] aes128/key[49] aes128/key[4] aes128/key[50] aes128/key[51]
+ aes128/key[52] aes128/key[53] aes128/key[54] aes128/key[55] aes128/key[56] aes128/key[57]
+ aes128/key[58] aes128/key[59] aes128/key[5] aes128/key[60] aes128/key[61] aes128/key[62]
+ aes128/key[63] aes128/key[64] aes128/key[65] aes128/key[66] aes128/key[67] aes128/key[68]
+ aes128/key[69] aes128/key[6] aes128/key[70] aes128/key[71] aes128/key[72] aes128/key[73]
+ aes128/key[74] aes128/key[75] aes128/key[76] aes128/key[77] aes128/key[78] aes128/key[79]
+ aes128/key[7] aes128/key[80] aes128/key[81] aes128/key[82] aes128/key[83] aes128/key[84]
+ aes128/key[85] aes128/key[86] aes128/key[87] aes128/key[88] aes128/key[89] aes128/key[8]
+ aes128/key[90] aes128/key[91] aes128/key[92] aes128/key[93] aes128/key[94] aes128/key[95]
+ aes128/key[96] aes128/key[97] aes128/key[98] aes128/key[99] aes128/key[9] aes128/out[0]
+ aes128/out[100] aes128/out[101] aes128/out[102] aes128/out[103] aes128/out[104]
+ aes128/out[105] aes128/out[106] aes128/out[107] aes128/out[108] aes128/out[109]
+ aes128/out[10] aes128/out[110] aes128/out[111] aes128/out[112] aes128/out[113] aes128/out[114]
+ aes128/out[115] aes128/out[116] aes128/out[117] aes128/out[118] aes128/out[119]
+ aes128/out[11] aes128/out[120] aes128/out[121] aes128/out[122] aes128/out[123] aes128/out[124]
+ aes128/out[125] aes128/out[126] aes128/out[127] aes128/out[12] aes128/out[13] aes128/out[14]
+ aes128/out[15] aes128/out[16] aes128/out[17] aes128/out[18] aes128/out[19] aes128/out[1]
+ aes128/out[20] aes128/out[21] aes128/out[22] aes128/out[23] aes128/out[24] aes128/out[25]
+ aes128/out[26] aes128/out[27] aes128/out[28] aes128/out[29] aes128/out[2] aes128/out[30]
+ aes128/out[31] aes128/out[32] aes128/out[33] aes128/out[34] aes128/out[35] aes128/out[36]
+ aes128/out[37] aes128/out[38] aes128/out[39] aes128/out[3] aes128/out[40] aes128/out[41]
+ aes128/out[42] aes128/out[43] aes128/out[44] aes128/out[45] aes128/out[46] aes128/out[47]
+ aes128/out[48] aes128/out[49] aes128/out[4] aes128/out[50] aes128/out[51] aes128/out[52]
+ aes128/out[53] aes128/out[54] aes128/out[55] aes128/out[56] aes128/out[57] aes128/out[58]
+ aes128/out[59] aes128/out[5] aes128/out[60] aes128/out[61] aes128/out[62] aes128/out[63]
+ aes128/out[64] aes128/out[65] aes128/out[66] aes128/out[67] aes128/out[68] aes128/out[69]
+ aes128/out[6] aes128/out[70] aes128/out[71] aes128/out[72] aes128/out[73] aes128/out[74]
+ aes128/out[75] aes128/out[76] aes128/out[77] aes128/out[78] aes128/out[79] aes128/out[7]
+ aes128/out[80] aes128/out[81] aes128/out[82] aes128/out[83] aes128/out[84] aes128/out[85]
+ aes128/out[86] aes128/out[87] aes128/out[88] aes128/out[89] aes128/out[8] aes128/out[90]
+ aes128/out[91] aes128/out[92] aes128/out[93] aes128/out[94] aes128/out[95] aes128/out[96]
+ aes128/out[97] aes128/out[98] aes128/out[99] aes128/out[9] aes128/state[0] aes128/state[100]
+ aes128/state[101] aes128/state[102] aes128/state[103] aes128/state[104] aes128/state[105]
+ aes128/state[106] aes128/state[107] aes128/state[108] aes128/state[109] aes128/state[10]
+ aes128/state[110] aes128/state[111] aes128/state[112] aes128/state[113] aes128/state[114]
+ aes128/state[115] aes128/state[116] aes128/state[117] aes128/state[118] aes128/state[119]
+ aes128/state[11] aes128/state[120] aes128/state[121] aes128/state[122] aes128/state[123]
+ aes128/state[124] aes128/state[125] aes128/state[126] aes128/state[127] aes128/state[12]
+ aes128/state[13] aes128/state[14] aes128/state[15] aes128/state[16] aes128/state[17]
+ aes128/state[18] aes128/state[19] aes128/state[1] aes128/state[20] aes128/state[21]
+ aes128/state[22] aes128/state[23] aes128/state[24] aes128/state[25] aes128/state[26]
+ aes128/state[27] aes128/state[28] aes128/state[29] aes128/state[2] aes128/state[30]
+ aes128/state[31] aes128/state[32] aes128/state[33] aes128/state[34] aes128/state[35]
+ aes128/state[36] aes128/state[37] aes128/state[38] aes128/state[39] aes128/state[3]
+ aes128/state[40] aes128/state[41] aes128/state[42] aes128/state[43] aes128/state[44]
+ aes128/state[45] aes128/state[46] aes128/state[47] aes128/state[48] aes128/state[49]
+ aes128/state[4] aes128/state[50] aes128/state[51] aes128/state[52] aes128/state[53]
+ aes128/state[54] aes128/state[55] aes128/state[56] aes128/state[57] aes128/state[58]
+ aes128/state[59] aes128/state[5] aes128/state[60] aes128/state[61] aes128/state[62]
+ aes128/state[63] aes128/state[64] aes128/state[65] aes128/state[66] aes128/state[67]
+ aes128/state[68] aes128/state[69] aes128/state[6] aes128/state[70] aes128/state[71]
+ aes128/state[72] aes128/state[73] aes128/state[74] aes128/state[75] aes128/state[76]
+ aes128/state[77] aes128/state[78] aes128/state[79] aes128/state[7] aes128/state[80]
+ aes128/state[81] aes128/state[82] aes128/state[83] aes128/state[84] aes128/state[85]
+ aes128/state[86] aes128/state[87] aes128/state[88] aes128/state[89] aes128/state[8]
+ aes128/state[90] aes128/state[91] aes128/state[92] aes128/state[93] aes128/state[94]
+ aes128/state[95] aes128/state[96] aes128/state[97] aes128/state[98] aes128/state[99]
+ aes128/state[9] vdd vss aes128
.ends

