magic
tech gf180mcuC
magscale 1 10
timestamp 1670228407
<< metal2 >>
rect 11032 595560 11256 597000
rect 33096 595560 33320 597000
rect 55160 595560 55384 597000
rect 77224 595560 77448 597000
rect 99288 595560 99512 597000
rect 121352 595560 121576 597000
rect 143416 595560 143640 597000
rect 165480 595560 165704 597000
rect 187544 595560 187768 597000
rect 209608 595560 209832 597000
rect 231672 595560 231896 597000
rect 253736 595560 253960 597000
rect 275800 595560 276024 597000
rect 297864 595560 298088 597000
rect 319928 595560 320152 597000
rect 341992 595560 342216 597000
rect 364056 595560 364280 597000
rect 386120 595560 386344 597000
rect 408184 595560 408408 597000
rect 430248 595560 430472 597000
rect 452312 595560 452536 597000
rect 474376 595560 474600 597000
rect 496440 595560 496664 597000
rect 518504 595560 518728 597000
rect 540568 595560 540792 597000
rect 562632 595560 562856 597000
rect 584696 595560 584920 597000
rect 47852 237748 47908 237758
rect 11564 4228 11620 4238
rect 11564 480 11620 4172
rect 47852 4228 47908 237692
rect 47852 4162 47908 4172
rect 11368 392 11620 480
rect 11368 -960 11592 392
rect 13272 -960 13496 480
rect 15176 -960 15400 480
rect 17080 -960 17304 480
rect 18984 -960 19208 480
rect 20888 -960 21112 480
rect 22792 -960 23016 480
rect 24696 -960 24920 480
rect 26600 -960 26824 480
rect 28504 -960 28728 480
rect 30408 -960 30632 480
rect 32312 -960 32536 480
rect 34216 -960 34440 480
rect 36120 -960 36344 480
rect 38024 -960 38248 480
rect 39928 -960 40152 480
rect 41832 -960 42056 480
rect 43736 -960 43960 480
rect 45640 -960 45864 480
rect 47544 -960 47768 480
rect 49448 -960 49672 480
rect 51352 -960 51576 480
rect 53256 -960 53480 480
rect 55160 -960 55384 480
rect 57064 -960 57288 480
rect 58968 -960 59192 480
rect 60872 -960 61096 480
rect 62776 -960 63000 480
rect 64680 -960 64904 480
rect 66584 -960 66808 480
rect 68488 -960 68712 480
rect 70392 -960 70616 480
rect 72296 -960 72520 480
rect 74200 -960 74424 480
rect 76104 -960 76328 480
rect 78008 -960 78232 480
rect 79912 -960 80136 480
rect 81816 -960 82040 480
rect 83720 -960 83944 480
rect 85624 -960 85848 480
rect 87528 -960 87752 480
rect 89432 -960 89656 480
rect 91336 -960 91560 480
rect 93240 -960 93464 480
rect 95144 -960 95368 480
rect 97048 -960 97272 480
rect 98952 -960 99176 480
rect 100856 -960 101080 480
rect 102760 -960 102984 480
rect 104664 -960 104888 480
rect 106568 -960 106792 480
rect 108472 -960 108696 480
rect 110376 -960 110600 480
rect 112280 -960 112504 480
rect 114184 -960 114408 480
rect 116088 -960 116312 480
rect 117992 -960 118216 480
rect 119896 -960 120120 480
rect 121800 -960 122024 480
rect 123704 -960 123928 480
rect 125608 -960 125832 480
rect 127512 -960 127736 480
rect 129416 -960 129640 480
rect 131320 -960 131544 480
rect 133224 -960 133448 480
rect 135128 -960 135352 480
rect 137032 -960 137256 480
rect 138936 -960 139160 480
rect 140840 -960 141064 480
rect 142744 -960 142968 480
rect 144648 -960 144872 480
rect 146552 -960 146776 480
rect 148456 -960 148680 480
rect 150360 -960 150584 480
rect 152264 -960 152488 480
rect 154168 -960 154392 480
rect 156072 -960 156296 480
rect 157976 -960 158200 480
rect 159880 -960 160104 480
rect 161784 -960 162008 480
rect 163688 -960 163912 480
rect 165592 -960 165816 480
rect 167496 -960 167720 480
rect 169400 -960 169624 480
rect 171304 -960 171528 480
rect 173208 -960 173432 480
rect 175112 -960 175336 480
rect 177016 -960 177240 480
rect 178920 -960 179144 480
rect 180824 -960 181048 480
rect 182728 -960 182952 480
rect 184632 -960 184856 480
rect 186536 -960 186760 480
rect 188440 -960 188664 480
rect 190344 -960 190568 480
rect 192248 -960 192472 480
rect 194152 -960 194376 480
rect 196056 -960 196280 480
rect 197960 -960 198184 480
rect 199864 -960 200088 480
rect 201768 -960 201992 480
rect 203672 -960 203896 480
rect 205576 -960 205800 480
rect 207480 -960 207704 480
rect 209384 -960 209608 480
rect 211288 -960 211512 480
rect 213192 -960 213416 480
rect 215096 -960 215320 480
rect 217000 -960 217224 480
rect 218904 -960 219128 480
rect 220808 -960 221032 480
rect 222712 -960 222936 480
rect 224616 -960 224840 480
rect 226520 -960 226744 480
rect 228424 -960 228648 480
rect 230328 -960 230552 480
rect 232232 -960 232456 480
rect 234136 -960 234360 480
rect 236040 -960 236264 480
rect 237944 -960 238168 480
rect 239848 -960 240072 480
rect 241752 -960 241976 480
rect 243656 -960 243880 480
rect 245560 -960 245784 480
rect 247464 -960 247688 480
rect 249368 -960 249592 480
rect 251272 -960 251496 480
rect 253176 -960 253400 480
rect 255080 -960 255304 480
rect 256984 -960 257208 480
rect 258888 -960 259112 480
rect 260792 -960 261016 480
rect 262696 -960 262920 480
rect 264600 -960 264824 480
rect 266504 -960 266728 480
rect 268408 -960 268632 480
rect 270312 -960 270536 480
rect 272216 -960 272440 480
rect 274120 -960 274344 480
rect 276024 -960 276248 480
rect 277928 -960 278152 480
rect 279832 -960 280056 480
rect 281736 -960 281960 480
rect 283640 -960 283864 480
rect 285544 -960 285768 480
rect 287448 -960 287672 480
rect 289352 -960 289576 480
rect 291256 -960 291480 480
rect 293160 -960 293384 480
rect 295064 -960 295288 480
rect 296968 -960 297192 480
rect 298872 -960 299096 480
rect 300776 -960 301000 480
rect 302680 -960 302904 480
rect 304584 -960 304808 480
rect 306488 -960 306712 480
rect 308392 -960 308616 480
rect 310296 -960 310520 480
rect 312200 -960 312424 480
rect 314104 -960 314328 480
rect 316008 -960 316232 480
rect 317912 -960 318136 480
rect 319816 -960 320040 480
rect 321720 -960 321944 480
rect 323624 -960 323848 480
rect 325528 -960 325752 480
rect 327432 -960 327656 480
rect 329336 -960 329560 480
rect 331240 -960 331464 480
rect 333144 -960 333368 480
rect 335048 -960 335272 480
rect 336952 -960 337176 480
rect 338856 -960 339080 480
rect 340760 -960 340984 480
rect 342664 -960 342888 480
rect 344568 -960 344792 480
rect 346472 -960 346696 480
rect 348376 -960 348600 480
rect 350280 -960 350504 480
rect 352184 -960 352408 480
rect 354088 -960 354312 480
rect 355992 -960 356216 480
rect 357896 -960 358120 480
rect 359800 -960 360024 480
rect 361704 -960 361928 480
rect 363608 -960 363832 480
rect 365512 -960 365736 480
rect 367416 -960 367640 480
rect 369320 -960 369544 480
rect 371224 -960 371448 480
rect 373128 -960 373352 480
rect 375032 -960 375256 480
rect 376936 -960 377160 480
rect 378840 -960 379064 480
rect 380744 -960 380968 480
rect 382648 -960 382872 480
rect 384552 -960 384776 480
rect 386456 -960 386680 480
rect 388360 -960 388584 480
rect 390264 -960 390488 480
rect 392168 -960 392392 480
rect 394072 -960 394296 480
rect 395976 -960 396200 480
rect 397880 -960 398104 480
rect 399784 -960 400008 480
rect 401688 -960 401912 480
rect 403592 -960 403816 480
rect 405496 -960 405720 480
rect 407400 -960 407624 480
rect 409304 -960 409528 480
rect 411208 -960 411432 480
rect 413112 -960 413336 480
rect 415016 -960 415240 480
rect 416920 -960 417144 480
rect 418824 -960 419048 480
rect 420728 -960 420952 480
rect 422632 -960 422856 480
rect 424536 -960 424760 480
rect 426440 -960 426664 480
rect 428344 -960 428568 480
rect 430248 -960 430472 480
rect 432152 -960 432376 480
rect 434056 -960 434280 480
rect 435960 -960 436184 480
rect 437864 -960 438088 480
rect 439768 -960 439992 480
rect 441672 -960 441896 480
rect 443576 -960 443800 480
rect 445480 -960 445704 480
rect 447384 -960 447608 480
rect 449288 -960 449512 480
rect 451192 -960 451416 480
rect 453096 -960 453320 480
rect 455000 -960 455224 480
rect 456904 -960 457128 480
rect 458808 -960 459032 480
rect 460712 -960 460936 480
rect 462616 -960 462840 480
rect 464520 -960 464744 480
rect 466424 -960 466648 480
rect 468328 -960 468552 480
rect 470232 -960 470456 480
rect 472136 -960 472360 480
rect 474040 -960 474264 480
rect 475944 -960 476168 480
rect 477848 -960 478072 480
rect 479752 -960 479976 480
rect 481656 -960 481880 480
rect 483560 -960 483784 480
rect 485464 -960 485688 480
rect 487368 -960 487592 480
rect 489272 -960 489496 480
rect 491176 -960 491400 480
rect 493080 -960 493304 480
rect 494984 -960 495208 480
rect 496888 -960 497112 480
rect 498792 -960 499016 480
rect 500696 -960 500920 480
rect 502600 -960 502824 480
rect 504504 -960 504728 480
rect 506408 -960 506632 480
rect 508312 -960 508536 480
rect 510216 -960 510440 480
rect 512120 -960 512344 480
rect 514024 -960 514248 480
rect 515928 -960 516152 480
rect 517832 -960 518056 480
rect 519736 -960 519960 480
rect 521640 -960 521864 480
rect 523544 -960 523768 480
rect 525448 -960 525672 480
rect 527352 -960 527576 480
rect 529256 -960 529480 480
rect 531160 -960 531384 480
rect 533064 -960 533288 480
rect 534968 -960 535192 480
rect 536872 -960 537096 480
rect 538776 -960 539000 480
rect 540680 -960 540904 480
rect 542584 -960 542808 480
rect 544488 -960 544712 480
rect 546392 -960 546616 480
rect 548296 -960 548520 480
rect 550200 -960 550424 480
rect 552104 -960 552328 480
rect 554008 -960 554232 480
rect 555912 -960 556136 480
rect 557816 -960 558040 480
rect 559720 -960 559944 480
rect 561624 -960 561848 480
rect 563528 -960 563752 480
rect 565432 -960 565656 480
rect 567336 -960 567560 480
rect 569240 -960 569464 480
rect 571144 -960 571368 480
rect 573048 -960 573272 480
rect 574952 -960 575176 480
rect 576856 -960 577080 480
rect 578760 -960 578984 480
rect 580664 -960 580888 480
rect 582568 -960 582792 480
rect 584472 -960 584696 480
<< via2 >>
rect 47852 237692 47908 237748
rect 11564 4172 11620 4228
rect 47852 4172 47908 4228
<< metal3 >>
rect 595560 588616 597000 588840
rect -960 587160 480 587384
rect 595560 575400 597000 575624
rect -960 573048 480 573272
rect 595560 562184 597000 562408
rect -960 558936 480 559160
rect 595560 548968 597000 549192
rect -960 544824 480 545048
rect 595560 535752 597000 535976
rect -960 530712 480 530936
rect 595560 522536 597000 522760
rect -960 516600 480 516824
rect 595560 509320 597000 509544
rect -960 502488 480 502712
rect 595560 496104 597000 496328
rect -960 488376 480 488600
rect 595560 482888 597000 483112
rect -960 474264 480 474488
rect 595560 469672 597000 469896
rect -960 460152 480 460376
rect 595560 456456 597000 456680
rect -960 446040 480 446264
rect 595560 443240 597000 443464
rect -960 431928 480 432152
rect 595560 430024 597000 430248
rect -960 417816 480 418040
rect 595560 416808 597000 417032
rect -960 403704 480 403928
rect 595560 403592 597000 403816
rect 595560 390376 597000 390600
rect -960 389592 480 389816
rect 595560 377160 597000 377384
rect -960 375480 480 375704
rect 595560 363944 597000 364168
rect -960 361368 480 361592
rect 595560 350728 597000 350952
rect -960 347256 480 347480
rect 595560 337512 597000 337736
rect -960 333144 480 333368
rect 595560 324296 597000 324520
rect -960 319032 480 319256
rect 595560 311080 597000 311304
rect -960 304920 480 305144
rect 595560 297864 597000 298088
rect -960 290808 480 291032
rect 595560 284648 597000 284872
rect -960 276696 480 276920
rect 595560 271432 597000 271656
rect -960 262584 480 262808
rect 595560 258216 597000 258440
rect -960 248472 480 248696
rect 595560 245000 597000 245224
rect 50204 237748 50260 237758
rect 47842 237692 47852 237748
rect 47908 237692 49868 237748
rect 49924 237692 49934 237748
rect 50204 237682 50260 237692
rect -960 234360 480 234584
rect 595560 231784 597000 232008
rect -960 220248 480 220472
rect 595560 218568 597000 218792
rect -960 206136 480 206360
rect 595560 205352 597000 205576
rect -960 192024 480 192248
rect 595560 192136 597000 192360
rect 595560 178920 597000 179144
rect -960 177912 480 178136
rect 595560 165704 597000 165928
rect -960 163800 480 164024
rect 595560 152488 597000 152712
rect -960 149688 480 149912
rect 595560 139272 597000 139496
rect -960 135576 480 135800
rect 595560 126056 597000 126280
rect -960 121464 480 121688
rect 595560 112840 597000 113064
rect -960 107352 480 107576
rect 595560 99624 597000 99848
rect -960 93240 480 93464
rect 595560 86408 597000 86632
rect -960 79128 480 79352
rect 595560 73192 597000 73416
rect -960 65016 480 65240
rect 595560 59976 597000 60200
rect -960 50904 480 51128
rect 595560 46760 597000 46984
rect -960 36792 480 37016
rect 595560 33544 597000 33768
rect -960 22680 480 22904
rect 595560 20328 597000 20552
rect -960 8568 480 8792
rect 595560 7112 597000 7336
rect 11554 4172 11564 4228
rect 11620 4172 47852 4228
rect 47908 4172 47918 4228
<< via3 >>
rect 49868 237692 49924 237748
rect 50204 237692 50260 237748
<< metal4 >>
rect -1916 598172 -1296 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 -1296 598172
rect -1916 598048 -1296 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 -1296 598048
rect -1916 597924 -1296 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 -1296 597924
rect -1916 597800 -1296 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 -1296 597800
rect -1916 586350 -1296 597744
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 -1296 586350
rect -1916 586226 -1296 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 -1296 586226
rect -1916 586102 -1296 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 -1296 586102
rect -1916 585978 -1296 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 -1296 585978
rect -1916 568350 -1296 585922
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 -1296 568350
rect -1916 568226 -1296 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 -1296 568226
rect -1916 568102 -1296 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 -1296 568102
rect -1916 567978 -1296 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 -1296 567978
rect -1916 550350 -1296 567922
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 -1296 550350
rect -1916 550226 -1296 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 -1296 550226
rect -1916 550102 -1296 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 -1296 550102
rect -1916 549978 -1296 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 -1296 549978
rect -1916 532350 -1296 549922
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 -1296 532350
rect -1916 532226 -1296 532294
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 -1296 532226
rect -1916 532102 -1296 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 -1296 532102
rect -1916 531978 -1296 532046
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 -1296 531978
rect -1916 514350 -1296 531922
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 -1296 514350
rect -1916 514226 -1296 514294
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 -1296 514226
rect -1916 514102 -1296 514170
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 -1296 514102
rect -1916 513978 -1296 514046
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 -1296 513978
rect -1916 496350 -1296 513922
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 -1296 496350
rect -1916 496226 -1296 496294
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 -1296 496226
rect -1916 496102 -1296 496170
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 -1296 496102
rect -1916 495978 -1296 496046
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 -1296 495978
rect -1916 478350 -1296 495922
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 -1296 478350
rect -1916 478226 -1296 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 -1296 478226
rect -1916 478102 -1296 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 -1296 478102
rect -1916 477978 -1296 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 -1296 477978
rect -1916 460350 -1296 477922
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 -1296 460350
rect -1916 460226 -1296 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 -1296 460226
rect -1916 460102 -1296 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 -1296 460102
rect -1916 459978 -1296 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 -1296 459978
rect -1916 442350 -1296 459922
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 -1296 442350
rect -1916 442226 -1296 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 -1296 442226
rect -1916 442102 -1296 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 -1296 442102
rect -1916 441978 -1296 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 -1296 441978
rect -1916 424350 -1296 441922
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 -1296 424350
rect -1916 424226 -1296 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 -1296 424226
rect -1916 424102 -1296 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 -1296 424102
rect -1916 423978 -1296 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 -1296 423978
rect -1916 406350 -1296 423922
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 -1296 406350
rect -1916 406226 -1296 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 -1296 406226
rect -1916 406102 -1296 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 -1296 406102
rect -1916 405978 -1296 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 -1296 405978
rect -1916 388350 -1296 405922
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 -1296 388350
rect -1916 388226 -1296 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 -1296 388226
rect -1916 388102 -1296 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 -1296 388102
rect -1916 387978 -1296 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 -1296 387978
rect -1916 370350 -1296 387922
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 -1296 370350
rect -1916 370226 -1296 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 -1296 370226
rect -1916 370102 -1296 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 -1296 370102
rect -1916 369978 -1296 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 -1296 369978
rect -1916 352350 -1296 369922
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 -1296 352350
rect -1916 352226 -1296 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 -1296 352226
rect -1916 352102 -1296 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 -1296 352102
rect -1916 351978 -1296 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 -1296 351978
rect -1916 334350 -1296 351922
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 -1296 334350
rect -1916 334226 -1296 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 -1296 334226
rect -1916 334102 -1296 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 -1296 334102
rect -1916 333978 -1296 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 -1296 333978
rect -1916 316350 -1296 333922
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 -1296 316350
rect -1916 316226 -1296 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 -1296 316226
rect -1916 316102 -1296 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 -1296 316102
rect -1916 315978 -1296 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 -1296 315978
rect -1916 298350 -1296 315922
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 -1296 298350
rect -1916 298226 -1296 298294
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 -1296 298226
rect -1916 298102 -1296 298170
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 -1296 298102
rect -1916 297978 -1296 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 -1296 297978
rect -1916 280350 -1296 297922
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 -1296 280350
rect -1916 280226 -1296 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 -1296 280226
rect -1916 280102 -1296 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 -1296 280102
rect -1916 279978 -1296 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 -1296 279978
rect -1916 262350 -1296 279922
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 -1296 262350
rect -1916 262226 -1296 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 -1296 262226
rect -1916 262102 -1296 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 -1296 262102
rect -1916 261978 -1296 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 -1296 261978
rect -1916 244350 -1296 261922
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 -1296 244350
rect -1916 244226 -1296 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 -1296 244226
rect -1916 244102 -1296 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 -1296 244102
rect -1916 243978 -1296 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 -1296 243978
rect -1916 226350 -1296 243922
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 -1296 226350
rect -1916 226226 -1296 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 -1296 226226
rect -1916 226102 -1296 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 -1296 226102
rect -1916 225978 -1296 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 -1296 225978
rect -1916 208350 -1296 225922
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 -1296 208350
rect -1916 208226 -1296 208294
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 -1296 208226
rect -1916 208102 -1296 208170
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 -1296 208102
rect -1916 207978 -1296 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 -1296 207978
rect -1916 190350 -1296 207922
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 -1296 190350
rect -1916 190226 -1296 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 -1296 190226
rect -1916 190102 -1296 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 -1296 190102
rect -1916 189978 -1296 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 -1296 189978
rect -1916 172350 -1296 189922
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 -1296 172350
rect -1916 172226 -1296 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 -1296 172226
rect -1916 172102 -1296 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 -1296 172102
rect -1916 171978 -1296 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 -1296 171978
rect -1916 154350 -1296 171922
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 -1296 154350
rect -1916 154226 -1296 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 -1296 154226
rect -1916 154102 -1296 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 -1296 154102
rect -1916 153978 -1296 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 -1296 153978
rect -1916 136350 -1296 153922
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 -1296 136350
rect -1916 136226 -1296 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 -1296 136226
rect -1916 136102 -1296 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 -1296 136102
rect -1916 135978 -1296 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 -1296 135978
rect -1916 118350 -1296 135922
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 -1296 118350
rect -1916 118226 -1296 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 -1296 118226
rect -1916 118102 -1296 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 -1296 118102
rect -1916 117978 -1296 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 -1296 117978
rect -1916 100350 -1296 117922
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 -1296 100350
rect -1916 100226 -1296 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 -1296 100226
rect -1916 100102 -1296 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 -1296 100102
rect -1916 99978 -1296 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 -1296 99978
rect -1916 82350 -1296 99922
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 -1296 82350
rect -1916 82226 -1296 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 -1296 82226
rect -1916 82102 -1296 82170
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 -1296 82102
rect -1916 81978 -1296 82046
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 -1296 81978
rect -1916 64350 -1296 81922
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 -1296 64350
rect -1916 64226 -1296 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 -1296 64226
rect -1916 64102 -1296 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 -1296 64102
rect -1916 63978 -1296 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 -1296 63978
rect -1916 46350 -1296 63922
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 -1296 46350
rect -1916 46226 -1296 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 -1296 46226
rect -1916 46102 -1296 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 -1296 46102
rect -1916 45978 -1296 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 -1296 45978
rect -1916 28350 -1296 45922
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 -1296 28350
rect -1916 28226 -1296 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 -1296 28226
rect -1916 28102 -1296 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 -1296 28102
rect -1916 27978 -1296 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 -1296 27978
rect -1916 10350 -1296 27922
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 -1296 10350
rect -1916 10226 -1296 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 -1296 10226
rect -1916 10102 -1296 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 -1296 10102
rect -1916 9978 -1296 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 -1296 9978
rect -1916 -1120 -1296 9922
rect -956 597212 -336 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 -336 597212
rect -956 597088 -336 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 -336 597088
rect -956 596964 -336 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 -336 596964
rect -956 596840 -336 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 -336 596840
rect -956 580350 -336 596784
rect -956 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 -336 580350
rect -956 580226 -336 580294
rect -956 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 -336 580226
rect -956 580102 -336 580170
rect -956 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 -336 580102
rect -956 579978 -336 580046
rect -956 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 -336 579978
rect -956 562350 -336 579922
rect -956 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 -336 562350
rect -956 562226 -336 562294
rect -956 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 -336 562226
rect -956 562102 -336 562170
rect -956 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 -336 562102
rect -956 561978 -336 562046
rect -956 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 -336 561978
rect -956 544350 -336 561922
rect -956 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 -336 544350
rect -956 544226 -336 544294
rect -956 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 -336 544226
rect -956 544102 -336 544170
rect -956 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 -336 544102
rect -956 543978 -336 544046
rect -956 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 -336 543978
rect -956 526350 -336 543922
rect -956 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 -336 526350
rect -956 526226 -336 526294
rect -956 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 -336 526226
rect -956 526102 -336 526170
rect -956 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 -336 526102
rect -956 525978 -336 526046
rect -956 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 -336 525978
rect -956 508350 -336 525922
rect -956 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 -336 508350
rect -956 508226 -336 508294
rect -956 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 -336 508226
rect -956 508102 -336 508170
rect -956 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 -336 508102
rect -956 507978 -336 508046
rect -956 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 -336 507978
rect -956 490350 -336 507922
rect -956 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 -336 490350
rect -956 490226 -336 490294
rect -956 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 -336 490226
rect -956 490102 -336 490170
rect -956 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 -336 490102
rect -956 489978 -336 490046
rect -956 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 -336 489978
rect -956 472350 -336 489922
rect -956 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 -336 472350
rect -956 472226 -336 472294
rect -956 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 -336 472226
rect -956 472102 -336 472170
rect -956 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 -336 472102
rect -956 471978 -336 472046
rect -956 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 -336 471978
rect -956 454350 -336 471922
rect -956 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 -336 454350
rect -956 454226 -336 454294
rect -956 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 -336 454226
rect -956 454102 -336 454170
rect -956 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 -336 454102
rect -956 453978 -336 454046
rect -956 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 -336 453978
rect -956 436350 -336 453922
rect -956 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 -336 436350
rect -956 436226 -336 436294
rect -956 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 -336 436226
rect -956 436102 -336 436170
rect -956 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 -336 436102
rect -956 435978 -336 436046
rect -956 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 -336 435978
rect -956 418350 -336 435922
rect -956 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 -336 418350
rect -956 418226 -336 418294
rect -956 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 -336 418226
rect -956 418102 -336 418170
rect -956 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 -336 418102
rect -956 417978 -336 418046
rect -956 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 -336 417978
rect -956 400350 -336 417922
rect -956 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 -336 400350
rect -956 400226 -336 400294
rect -956 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 -336 400226
rect -956 400102 -336 400170
rect -956 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 -336 400102
rect -956 399978 -336 400046
rect -956 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 -336 399978
rect -956 382350 -336 399922
rect -956 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 -336 382350
rect -956 382226 -336 382294
rect -956 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 -336 382226
rect -956 382102 -336 382170
rect -956 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 -336 382102
rect -956 381978 -336 382046
rect -956 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 -336 381978
rect -956 364350 -336 381922
rect -956 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 -336 364350
rect -956 364226 -336 364294
rect -956 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 -336 364226
rect -956 364102 -336 364170
rect -956 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 -336 364102
rect -956 363978 -336 364046
rect -956 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 -336 363978
rect -956 346350 -336 363922
rect -956 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 -336 346350
rect -956 346226 -336 346294
rect -956 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 -336 346226
rect -956 346102 -336 346170
rect -956 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 -336 346102
rect -956 345978 -336 346046
rect -956 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 -336 345978
rect -956 328350 -336 345922
rect -956 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 -336 328350
rect -956 328226 -336 328294
rect -956 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 -336 328226
rect -956 328102 -336 328170
rect -956 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 -336 328102
rect -956 327978 -336 328046
rect -956 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 -336 327978
rect -956 310350 -336 327922
rect -956 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 -336 310350
rect -956 310226 -336 310294
rect -956 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 -336 310226
rect -956 310102 -336 310170
rect -956 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 -336 310102
rect -956 309978 -336 310046
rect -956 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 -336 309978
rect -956 292350 -336 309922
rect -956 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 -336 292350
rect -956 292226 -336 292294
rect -956 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 -336 292226
rect -956 292102 -336 292170
rect -956 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 -336 292102
rect -956 291978 -336 292046
rect -956 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 -336 291978
rect -956 274350 -336 291922
rect -956 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 -336 274350
rect -956 274226 -336 274294
rect -956 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 -336 274226
rect -956 274102 -336 274170
rect -956 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 -336 274102
rect -956 273978 -336 274046
rect -956 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 -336 273978
rect -956 256350 -336 273922
rect -956 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 -336 256350
rect -956 256226 -336 256294
rect -956 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 -336 256226
rect -956 256102 -336 256170
rect -956 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 -336 256102
rect -956 255978 -336 256046
rect -956 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 -336 255978
rect -956 238350 -336 255922
rect -956 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 -336 238350
rect -956 238226 -336 238294
rect -956 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 -336 238226
rect -956 238102 -336 238170
rect -956 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 -336 238102
rect -956 237978 -336 238046
rect -956 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 -336 237978
rect -956 220350 -336 237922
rect -956 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 -336 220350
rect -956 220226 -336 220294
rect -956 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 -336 220226
rect -956 220102 -336 220170
rect -956 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 -336 220102
rect -956 219978 -336 220046
rect -956 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 -336 219978
rect -956 202350 -336 219922
rect -956 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 -336 202350
rect -956 202226 -336 202294
rect -956 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 -336 202226
rect -956 202102 -336 202170
rect -956 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 -336 202102
rect -956 201978 -336 202046
rect -956 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 -336 201978
rect -956 184350 -336 201922
rect -956 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 -336 184350
rect -956 184226 -336 184294
rect -956 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 -336 184226
rect -956 184102 -336 184170
rect -956 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 -336 184102
rect -956 183978 -336 184046
rect -956 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 -336 183978
rect -956 166350 -336 183922
rect -956 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 -336 166350
rect -956 166226 -336 166294
rect -956 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 -336 166226
rect -956 166102 -336 166170
rect -956 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 -336 166102
rect -956 165978 -336 166046
rect -956 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 -336 165978
rect -956 148350 -336 165922
rect -956 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 -336 148350
rect -956 148226 -336 148294
rect -956 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 -336 148226
rect -956 148102 -336 148170
rect -956 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 -336 148102
rect -956 147978 -336 148046
rect -956 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 -336 147978
rect -956 130350 -336 147922
rect -956 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 -336 130350
rect -956 130226 -336 130294
rect -956 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 -336 130226
rect -956 130102 -336 130170
rect -956 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 -336 130102
rect -956 129978 -336 130046
rect -956 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 -336 129978
rect -956 112350 -336 129922
rect -956 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 -336 112350
rect -956 112226 -336 112294
rect -956 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 -336 112226
rect -956 112102 -336 112170
rect -956 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 -336 112102
rect -956 111978 -336 112046
rect -956 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 -336 111978
rect -956 94350 -336 111922
rect -956 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 -336 94350
rect -956 94226 -336 94294
rect -956 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 -336 94226
rect -956 94102 -336 94170
rect -956 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 -336 94102
rect -956 93978 -336 94046
rect -956 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 -336 93978
rect -956 76350 -336 93922
rect -956 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 -336 76350
rect -956 76226 -336 76294
rect -956 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 -336 76226
rect -956 76102 -336 76170
rect -956 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 -336 76102
rect -956 75978 -336 76046
rect -956 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 -336 75978
rect -956 58350 -336 75922
rect -956 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 -336 58350
rect -956 58226 -336 58294
rect -956 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 -336 58226
rect -956 58102 -336 58170
rect -956 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 -336 58102
rect -956 57978 -336 58046
rect -956 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 -336 57978
rect -956 40350 -336 57922
rect -956 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 -336 40350
rect -956 40226 -336 40294
rect -956 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 -336 40226
rect -956 40102 -336 40170
rect -956 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 -336 40102
rect -956 39978 -336 40046
rect -956 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 -336 39978
rect -956 22350 -336 39922
rect -956 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 -336 22350
rect -956 22226 -336 22294
rect -956 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 -336 22226
rect -956 22102 -336 22170
rect -956 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 -336 22102
rect -956 21978 -336 22046
rect -956 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 -336 21978
rect -956 4350 -336 21922
rect -956 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 -336 4350
rect -956 4226 -336 4294
rect -956 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 -336 4226
rect -956 4102 -336 4170
rect -956 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 -336 4102
rect -956 3978 -336 4046
rect -956 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 -336 3978
rect -956 -160 -336 3922
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 -336 -160
rect -956 -284 -336 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 -336 -284
rect -956 -408 -336 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 -336 -408
rect -956 -532 -336 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 -336 -532
rect -956 -684 -336 -588
rect 3154 597212 3774 598268
rect 3154 597156 3250 597212
rect 3306 597156 3374 597212
rect 3430 597156 3498 597212
rect 3554 597156 3622 597212
rect 3678 597156 3774 597212
rect 3154 597088 3774 597156
rect 3154 597032 3250 597088
rect 3306 597032 3374 597088
rect 3430 597032 3498 597088
rect 3554 597032 3622 597088
rect 3678 597032 3774 597088
rect 3154 596964 3774 597032
rect 3154 596908 3250 596964
rect 3306 596908 3374 596964
rect 3430 596908 3498 596964
rect 3554 596908 3622 596964
rect 3678 596908 3774 596964
rect 3154 596840 3774 596908
rect 3154 596784 3250 596840
rect 3306 596784 3374 596840
rect 3430 596784 3498 596840
rect 3554 596784 3622 596840
rect 3678 596784 3774 596840
rect 3154 580350 3774 596784
rect 3154 580294 3250 580350
rect 3306 580294 3374 580350
rect 3430 580294 3498 580350
rect 3554 580294 3622 580350
rect 3678 580294 3774 580350
rect 3154 580226 3774 580294
rect 3154 580170 3250 580226
rect 3306 580170 3374 580226
rect 3430 580170 3498 580226
rect 3554 580170 3622 580226
rect 3678 580170 3774 580226
rect 3154 580102 3774 580170
rect 3154 580046 3250 580102
rect 3306 580046 3374 580102
rect 3430 580046 3498 580102
rect 3554 580046 3622 580102
rect 3678 580046 3774 580102
rect 3154 579978 3774 580046
rect 3154 579922 3250 579978
rect 3306 579922 3374 579978
rect 3430 579922 3498 579978
rect 3554 579922 3622 579978
rect 3678 579922 3774 579978
rect 3154 562350 3774 579922
rect 3154 562294 3250 562350
rect 3306 562294 3374 562350
rect 3430 562294 3498 562350
rect 3554 562294 3622 562350
rect 3678 562294 3774 562350
rect 3154 562226 3774 562294
rect 3154 562170 3250 562226
rect 3306 562170 3374 562226
rect 3430 562170 3498 562226
rect 3554 562170 3622 562226
rect 3678 562170 3774 562226
rect 3154 562102 3774 562170
rect 3154 562046 3250 562102
rect 3306 562046 3374 562102
rect 3430 562046 3498 562102
rect 3554 562046 3622 562102
rect 3678 562046 3774 562102
rect 3154 561978 3774 562046
rect 3154 561922 3250 561978
rect 3306 561922 3374 561978
rect 3430 561922 3498 561978
rect 3554 561922 3622 561978
rect 3678 561922 3774 561978
rect 3154 544350 3774 561922
rect 3154 544294 3250 544350
rect 3306 544294 3374 544350
rect 3430 544294 3498 544350
rect 3554 544294 3622 544350
rect 3678 544294 3774 544350
rect 3154 544226 3774 544294
rect 3154 544170 3250 544226
rect 3306 544170 3374 544226
rect 3430 544170 3498 544226
rect 3554 544170 3622 544226
rect 3678 544170 3774 544226
rect 3154 544102 3774 544170
rect 3154 544046 3250 544102
rect 3306 544046 3374 544102
rect 3430 544046 3498 544102
rect 3554 544046 3622 544102
rect 3678 544046 3774 544102
rect 3154 543978 3774 544046
rect 3154 543922 3250 543978
rect 3306 543922 3374 543978
rect 3430 543922 3498 543978
rect 3554 543922 3622 543978
rect 3678 543922 3774 543978
rect 3154 526350 3774 543922
rect 3154 526294 3250 526350
rect 3306 526294 3374 526350
rect 3430 526294 3498 526350
rect 3554 526294 3622 526350
rect 3678 526294 3774 526350
rect 3154 526226 3774 526294
rect 3154 526170 3250 526226
rect 3306 526170 3374 526226
rect 3430 526170 3498 526226
rect 3554 526170 3622 526226
rect 3678 526170 3774 526226
rect 3154 526102 3774 526170
rect 3154 526046 3250 526102
rect 3306 526046 3374 526102
rect 3430 526046 3498 526102
rect 3554 526046 3622 526102
rect 3678 526046 3774 526102
rect 3154 525978 3774 526046
rect 3154 525922 3250 525978
rect 3306 525922 3374 525978
rect 3430 525922 3498 525978
rect 3554 525922 3622 525978
rect 3678 525922 3774 525978
rect 3154 508350 3774 525922
rect 3154 508294 3250 508350
rect 3306 508294 3374 508350
rect 3430 508294 3498 508350
rect 3554 508294 3622 508350
rect 3678 508294 3774 508350
rect 3154 508226 3774 508294
rect 3154 508170 3250 508226
rect 3306 508170 3374 508226
rect 3430 508170 3498 508226
rect 3554 508170 3622 508226
rect 3678 508170 3774 508226
rect 3154 508102 3774 508170
rect 3154 508046 3250 508102
rect 3306 508046 3374 508102
rect 3430 508046 3498 508102
rect 3554 508046 3622 508102
rect 3678 508046 3774 508102
rect 3154 507978 3774 508046
rect 3154 507922 3250 507978
rect 3306 507922 3374 507978
rect 3430 507922 3498 507978
rect 3554 507922 3622 507978
rect 3678 507922 3774 507978
rect 3154 490350 3774 507922
rect 3154 490294 3250 490350
rect 3306 490294 3374 490350
rect 3430 490294 3498 490350
rect 3554 490294 3622 490350
rect 3678 490294 3774 490350
rect 3154 490226 3774 490294
rect 3154 490170 3250 490226
rect 3306 490170 3374 490226
rect 3430 490170 3498 490226
rect 3554 490170 3622 490226
rect 3678 490170 3774 490226
rect 3154 490102 3774 490170
rect 3154 490046 3250 490102
rect 3306 490046 3374 490102
rect 3430 490046 3498 490102
rect 3554 490046 3622 490102
rect 3678 490046 3774 490102
rect 3154 489978 3774 490046
rect 3154 489922 3250 489978
rect 3306 489922 3374 489978
rect 3430 489922 3498 489978
rect 3554 489922 3622 489978
rect 3678 489922 3774 489978
rect 3154 472350 3774 489922
rect 3154 472294 3250 472350
rect 3306 472294 3374 472350
rect 3430 472294 3498 472350
rect 3554 472294 3622 472350
rect 3678 472294 3774 472350
rect 3154 472226 3774 472294
rect 3154 472170 3250 472226
rect 3306 472170 3374 472226
rect 3430 472170 3498 472226
rect 3554 472170 3622 472226
rect 3678 472170 3774 472226
rect 3154 472102 3774 472170
rect 3154 472046 3250 472102
rect 3306 472046 3374 472102
rect 3430 472046 3498 472102
rect 3554 472046 3622 472102
rect 3678 472046 3774 472102
rect 3154 471978 3774 472046
rect 3154 471922 3250 471978
rect 3306 471922 3374 471978
rect 3430 471922 3498 471978
rect 3554 471922 3622 471978
rect 3678 471922 3774 471978
rect 3154 454350 3774 471922
rect 3154 454294 3250 454350
rect 3306 454294 3374 454350
rect 3430 454294 3498 454350
rect 3554 454294 3622 454350
rect 3678 454294 3774 454350
rect 3154 454226 3774 454294
rect 3154 454170 3250 454226
rect 3306 454170 3374 454226
rect 3430 454170 3498 454226
rect 3554 454170 3622 454226
rect 3678 454170 3774 454226
rect 3154 454102 3774 454170
rect 3154 454046 3250 454102
rect 3306 454046 3374 454102
rect 3430 454046 3498 454102
rect 3554 454046 3622 454102
rect 3678 454046 3774 454102
rect 3154 453978 3774 454046
rect 3154 453922 3250 453978
rect 3306 453922 3374 453978
rect 3430 453922 3498 453978
rect 3554 453922 3622 453978
rect 3678 453922 3774 453978
rect 3154 436350 3774 453922
rect 3154 436294 3250 436350
rect 3306 436294 3374 436350
rect 3430 436294 3498 436350
rect 3554 436294 3622 436350
rect 3678 436294 3774 436350
rect 3154 436226 3774 436294
rect 3154 436170 3250 436226
rect 3306 436170 3374 436226
rect 3430 436170 3498 436226
rect 3554 436170 3622 436226
rect 3678 436170 3774 436226
rect 3154 436102 3774 436170
rect 3154 436046 3250 436102
rect 3306 436046 3374 436102
rect 3430 436046 3498 436102
rect 3554 436046 3622 436102
rect 3678 436046 3774 436102
rect 3154 435978 3774 436046
rect 3154 435922 3250 435978
rect 3306 435922 3374 435978
rect 3430 435922 3498 435978
rect 3554 435922 3622 435978
rect 3678 435922 3774 435978
rect 3154 418350 3774 435922
rect 3154 418294 3250 418350
rect 3306 418294 3374 418350
rect 3430 418294 3498 418350
rect 3554 418294 3622 418350
rect 3678 418294 3774 418350
rect 3154 418226 3774 418294
rect 3154 418170 3250 418226
rect 3306 418170 3374 418226
rect 3430 418170 3498 418226
rect 3554 418170 3622 418226
rect 3678 418170 3774 418226
rect 3154 418102 3774 418170
rect 3154 418046 3250 418102
rect 3306 418046 3374 418102
rect 3430 418046 3498 418102
rect 3554 418046 3622 418102
rect 3678 418046 3774 418102
rect 3154 417978 3774 418046
rect 3154 417922 3250 417978
rect 3306 417922 3374 417978
rect 3430 417922 3498 417978
rect 3554 417922 3622 417978
rect 3678 417922 3774 417978
rect 3154 400350 3774 417922
rect 3154 400294 3250 400350
rect 3306 400294 3374 400350
rect 3430 400294 3498 400350
rect 3554 400294 3622 400350
rect 3678 400294 3774 400350
rect 3154 400226 3774 400294
rect 3154 400170 3250 400226
rect 3306 400170 3374 400226
rect 3430 400170 3498 400226
rect 3554 400170 3622 400226
rect 3678 400170 3774 400226
rect 3154 400102 3774 400170
rect 3154 400046 3250 400102
rect 3306 400046 3374 400102
rect 3430 400046 3498 400102
rect 3554 400046 3622 400102
rect 3678 400046 3774 400102
rect 3154 399978 3774 400046
rect 3154 399922 3250 399978
rect 3306 399922 3374 399978
rect 3430 399922 3498 399978
rect 3554 399922 3622 399978
rect 3678 399922 3774 399978
rect 3154 382350 3774 399922
rect 3154 382294 3250 382350
rect 3306 382294 3374 382350
rect 3430 382294 3498 382350
rect 3554 382294 3622 382350
rect 3678 382294 3774 382350
rect 3154 382226 3774 382294
rect 3154 382170 3250 382226
rect 3306 382170 3374 382226
rect 3430 382170 3498 382226
rect 3554 382170 3622 382226
rect 3678 382170 3774 382226
rect 3154 382102 3774 382170
rect 3154 382046 3250 382102
rect 3306 382046 3374 382102
rect 3430 382046 3498 382102
rect 3554 382046 3622 382102
rect 3678 382046 3774 382102
rect 3154 381978 3774 382046
rect 3154 381922 3250 381978
rect 3306 381922 3374 381978
rect 3430 381922 3498 381978
rect 3554 381922 3622 381978
rect 3678 381922 3774 381978
rect 3154 364350 3774 381922
rect 3154 364294 3250 364350
rect 3306 364294 3374 364350
rect 3430 364294 3498 364350
rect 3554 364294 3622 364350
rect 3678 364294 3774 364350
rect 3154 364226 3774 364294
rect 3154 364170 3250 364226
rect 3306 364170 3374 364226
rect 3430 364170 3498 364226
rect 3554 364170 3622 364226
rect 3678 364170 3774 364226
rect 3154 364102 3774 364170
rect 3154 364046 3250 364102
rect 3306 364046 3374 364102
rect 3430 364046 3498 364102
rect 3554 364046 3622 364102
rect 3678 364046 3774 364102
rect 3154 363978 3774 364046
rect 3154 363922 3250 363978
rect 3306 363922 3374 363978
rect 3430 363922 3498 363978
rect 3554 363922 3622 363978
rect 3678 363922 3774 363978
rect 3154 346350 3774 363922
rect 3154 346294 3250 346350
rect 3306 346294 3374 346350
rect 3430 346294 3498 346350
rect 3554 346294 3622 346350
rect 3678 346294 3774 346350
rect 3154 346226 3774 346294
rect 3154 346170 3250 346226
rect 3306 346170 3374 346226
rect 3430 346170 3498 346226
rect 3554 346170 3622 346226
rect 3678 346170 3774 346226
rect 3154 346102 3774 346170
rect 3154 346046 3250 346102
rect 3306 346046 3374 346102
rect 3430 346046 3498 346102
rect 3554 346046 3622 346102
rect 3678 346046 3774 346102
rect 3154 345978 3774 346046
rect 3154 345922 3250 345978
rect 3306 345922 3374 345978
rect 3430 345922 3498 345978
rect 3554 345922 3622 345978
rect 3678 345922 3774 345978
rect 3154 328350 3774 345922
rect 3154 328294 3250 328350
rect 3306 328294 3374 328350
rect 3430 328294 3498 328350
rect 3554 328294 3622 328350
rect 3678 328294 3774 328350
rect 3154 328226 3774 328294
rect 3154 328170 3250 328226
rect 3306 328170 3374 328226
rect 3430 328170 3498 328226
rect 3554 328170 3622 328226
rect 3678 328170 3774 328226
rect 3154 328102 3774 328170
rect 3154 328046 3250 328102
rect 3306 328046 3374 328102
rect 3430 328046 3498 328102
rect 3554 328046 3622 328102
rect 3678 328046 3774 328102
rect 3154 327978 3774 328046
rect 3154 327922 3250 327978
rect 3306 327922 3374 327978
rect 3430 327922 3498 327978
rect 3554 327922 3622 327978
rect 3678 327922 3774 327978
rect 3154 310350 3774 327922
rect 3154 310294 3250 310350
rect 3306 310294 3374 310350
rect 3430 310294 3498 310350
rect 3554 310294 3622 310350
rect 3678 310294 3774 310350
rect 3154 310226 3774 310294
rect 3154 310170 3250 310226
rect 3306 310170 3374 310226
rect 3430 310170 3498 310226
rect 3554 310170 3622 310226
rect 3678 310170 3774 310226
rect 3154 310102 3774 310170
rect 3154 310046 3250 310102
rect 3306 310046 3374 310102
rect 3430 310046 3498 310102
rect 3554 310046 3622 310102
rect 3678 310046 3774 310102
rect 3154 309978 3774 310046
rect 3154 309922 3250 309978
rect 3306 309922 3374 309978
rect 3430 309922 3498 309978
rect 3554 309922 3622 309978
rect 3678 309922 3774 309978
rect 3154 292350 3774 309922
rect 3154 292294 3250 292350
rect 3306 292294 3374 292350
rect 3430 292294 3498 292350
rect 3554 292294 3622 292350
rect 3678 292294 3774 292350
rect 3154 292226 3774 292294
rect 3154 292170 3250 292226
rect 3306 292170 3374 292226
rect 3430 292170 3498 292226
rect 3554 292170 3622 292226
rect 3678 292170 3774 292226
rect 3154 292102 3774 292170
rect 3154 292046 3250 292102
rect 3306 292046 3374 292102
rect 3430 292046 3498 292102
rect 3554 292046 3622 292102
rect 3678 292046 3774 292102
rect 3154 291978 3774 292046
rect 3154 291922 3250 291978
rect 3306 291922 3374 291978
rect 3430 291922 3498 291978
rect 3554 291922 3622 291978
rect 3678 291922 3774 291978
rect 3154 274350 3774 291922
rect 3154 274294 3250 274350
rect 3306 274294 3374 274350
rect 3430 274294 3498 274350
rect 3554 274294 3622 274350
rect 3678 274294 3774 274350
rect 3154 274226 3774 274294
rect 3154 274170 3250 274226
rect 3306 274170 3374 274226
rect 3430 274170 3498 274226
rect 3554 274170 3622 274226
rect 3678 274170 3774 274226
rect 3154 274102 3774 274170
rect 3154 274046 3250 274102
rect 3306 274046 3374 274102
rect 3430 274046 3498 274102
rect 3554 274046 3622 274102
rect 3678 274046 3774 274102
rect 3154 273978 3774 274046
rect 3154 273922 3250 273978
rect 3306 273922 3374 273978
rect 3430 273922 3498 273978
rect 3554 273922 3622 273978
rect 3678 273922 3774 273978
rect 3154 256350 3774 273922
rect 3154 256294 3250 256350
rect 3306 256294 3374 256350
rect 3430 256294 3498 256350
rect 3554 256294 3622 256350
rect 3678 256294 3774 256350
rect 3154 256226 3774 256294
rect 3154 256170 3250 256226
rect 3306 256170 3374 256226
rect 3430 256170 3498 256226
rect 3554 256170 3622 256226
rect 3678 256170 3774 256226
rect 3154 256102 3774 256170
rect 3154 256046 3250 256102
rect 3306 256046 3374 256102
rect 3430 256046 3498 256102
rect 3554 256046 3622 256102
rect 3678 256046 3774 256102
rect 3154 255978 3774 256046
rect 3154 255922 3250 255978
rect 3306 255922 3374 255978
rect 3430 255922 3498 255978
rect 3554 255922 3622 255978
rect 3678 255922 3774 255978
rect 3154 238350 3774 255922
rect 3154 238294 3250 238350
rect 3306 238294 3374 238350
rect 3430 238294 3498 238350
rect 3554 238294 3622 238350
rect 3678 238294 3774 238350
rect 3154 238226 3774 238294
rect 3154 238170 3250 238226
rect 3306 238170 3374 238226
rect 3430 238170 3498 238226
rect 3554 238170 3622 238226
rect 3678 238170 3774 238226
rect 3154 238102 3774 238170
rect 3154 238046 3250 238102
rect 3306 238046 3374 238102
rect 3430 238046 3498 238102
rect 3554 238046 3622 238102
rect 3678 238046 3774 238102
rect 3154 237978 3774 238046
rect 3154 237922 3250 237978
rect 3306 237922 3374 237978
rect 3430 237922 3498 237978
rect 3554 237922 3622 237978
rect 3678 237922 3774 237978
rect 3154 220350 3774 237922
rect 3154 220294 3250 220350
rect 3306 220294 3374 220350
rect 3430 220294 3498 220350
rect 3554 220294 3622 220350
rect 3678 220294 3774 220350
rect 3154 220226 3774 220294
rect 3154 220170 3250 220226
rect 3306 220170 3374 220226
rect 3430 220170 3498 220226
rect 3554 220170 3622 220226
rect 3678 220170 3774 220226
rect 3154 220102 3774 220170
rect 3154 220046 3250 220102
rect 3306 220046 3374 220102
rect 3430 220046 3498 220102
rect 3554 220046 3622 220102
rect 3678 220046 3774 220102
rect 3154 219978 3774 220046
rect 3154 219922 3250 219978
rect 3306 219922 3374 219978
rect 3430 219922 3498 219978
rect 3554 219922 3622 219978
rect 3678 219922 3774 219978
rect 3154 202350 3774 219922
rect 3154 202294 3250 202350
rect 3306 202294 3374 202350
rect 3430 202294 3498 202350
rect 3554 202294 3622 202350
rect 3678 202294 3774 202350
rect 3154 202226 3774 202294
rect 3154 202170 3250 202226
rect 3306 202170 3374 202226
rect 3430 202170 3498 202226
rect 3554 202170 3622 202226
rect 3678 202170 3774 202226
rect 3154 202102 3774 202170
rect 3154 202046 3250 202102
rect 3306 202046 3374 202102
rect 3430 202046 3498 202102
rect 3554 202046 3622 202102
rect 3678 202046 3774 202102
rect 3154 201978 3774 202046
rect 3154 201922 3250 201978
rect 3306 201922 3374 201978
rect 3430 201922 3498 201978
rect 3554 201922 3622 201978
rect 3678 201922 3774 201978
rect 3154 184350 3774 201922
rect 3154 184294 3250 184350
rect 3306 184294 3374 184350
rect 3430 184294 3498 184350
rect 3554 184294 3622 184350
rect 3678 184294 3774 184350
rect 3154 184226 3774 184294
rect 3154 184170 3250 184226
rect 3306 184170 3374 184226
rect 3430 184170 3498 184226
rect 3554 184170 3622 184226
rect 3678 184170 3774 184226
rect 3154 184102 3774 184170
rect 3154 184046 3250 184102
rect 3306 184046 3374 184102
rect 3430 184046 3498 184102
rect 3554 184046 3622 184102
rect 3678 184046 3774 184102
rect 3154 183978 3774 184046
rect 3154 183922 3250 183978
rect 3306 183922 3374 183978
rect 3430 183922 3498 183978
rect 3554 183922 3622 183978
rect 3678 183922 3774 183978
rect 3154 166350 3774 183922
rect 3154 166294 3250 166350
rect 3306 166294 3374 166350
rect 3430 166294 3498 166350
rect 3554 166294 3622 166350
rect 3678 166294 3774 166350
rect 3154 166226 3774 166294
rect 3154 166170 3250 166226
rect 3306 166170 3374 166226
rect 3430 166170 3498 166226
rect 3554 166170 3622 166226
rect 3678 166170 3774 166226
rect 3154 166102 3774 166170
rect 3154 166046 3250 166102
rect 3306 166046 3374 166102
rect 3430 166046 3498 166102
rect 3554 166046 3622 166102
rect 3678 166046 3774 166102
rect 3154 165978 3774 166046
rect 3154 165922 3250 165978
rect 3306 165922 3374 165978
rect 3430 165922 3498 165978
rect 3554 165922 3622 165978
rect 3678 165922 3774 165978
rect 3154 148350 3774 165922
rect 3154 148294 3250 148350
rect 3306 148294 3374 148350
rect 3430 148294 3498 148350
rect 3554 148294 3622 148350
rect 3678 148294 3774 148350
rect 3154 148226 3774 148294
rect 3154 148170 3250 148226
rect 3306 148170 3374 148226
rect 3430 148170 3498 148226
rect 3554 148170 3622 148226
rect 3678 148170 3774 148226
rect 3154 148102 3774 148170
rect 3154 148046 3250 148102
rect 3306 148046 3374 148102
rect 3430 148046 3498 148102
rect 3554 148046 3622 148102
rect 3678 148046 3774 148102
rect 3154 147978 3774 148046
rect 3154 147922 3250 147978
rect 3306 147922 3374 147978
rect 3430 147922 3498 147978
rect 3554 147922 3622 147978
rect 3678 147922 3774 147978
rect 3154 130350 3774 147922
rect 3154 130294 3250 130350
rect 3306 130294 3374 130350
rect 3430 130294 3498 130350
rect 3554 130294 3622 130350
rect 3678 130294 3774 130350
rect 3154 130226 3774 130294
rect 3154 130170 3250 130226
rect 3306 130170 3374 130226
rect 3430 130170 3498 130226
rect 3554 130170 3622 130226
rect 3678 130170 3774 130226
rect 3154 130102 3774 130170
rect 3154 130046 3250 130102
rect 3306 130046 3374 130102
rect 3430 130046 3498 130102
rect 3554 130046 3622 130102
rect 3678 130046 3774 130102
rect 3154 129978 3774 130046
rect 3154 129922 3250 129978
rect 3306 129922 3374 129978
rect 3430 129922 3498 129978
rect 3554 129922 3622 129978
rect 3678 129922 3774 129978
rect 3154 112350 3774 129922
rect 3154 112294 3250 112350
rect 3306 112294 3374 112350
rect 3430 112294 3498 112350
rect 3554 112294 3622 112350
rect 3678 112294 3774 112350
rect 3154 112226 3774 112294
rect 3154 112170 3250 112226
rect 3306 112170 3374 112226
rect 3430 112170 3498 112226
rect 3554 112170 3622 112226
rect 3678 112170 3774 112226
rect 3154 112102 3774 112170
rect 3154 112046 3250 112102
rect 3306 112046 3374 112102
rect 3430 112046 3498 112102
rect 3554 112046 3622 112102
rect 3678 112046 3774 112102
rect 3154 111978 3774 112046
rect 3154 111922 3250 111978
rect 3306 111922 3374 111978
rect 3430 111922 3498 111978
rect 3554 111922 3622 111978
rect 3678 111922 3774 111978
rect 3154 94350 3774 111922
rect 3154 94294 3250 94350
rect 3306 94294 3374 94350
rect 3430 94294 3498 94350
rect 3554 94294 3622 94350
rect 3678 94294 3774 94350
rect 3154 94226 3774 94294
rect 3154 94170 3250 94226
rect 3306 94170 3374 94226
rect 3430 94170 3498 94226
rect 3554 94170 3622 94226
rect 3678 94170 3774 94226
rect 3154 94102 3774 94170
rect 3154 94046 3250 94102
rect 3306 94046 3374 94102
rect 3430 94046 3498 94102
rect 3554 94046 3622 94102
rect 3678 94046 3774 94102
rect 3154 93978 3774 94046
rect 3154 93922 3250 93978
rect 3306 93922 3374 93978
rect 3430 93922 3498 93978
rect 3554 93922 3622 93978
rect 3678 93922 3774 93978
rect 3154 76350 3774 93922
rect 3154 76294 3250 76350
rect 3306 76294 3374 76350
rect 3430 76294 3498 76350
rect 3554 76294 3622 76350
rect 3678 76294 3774 76350
rect 3154 76226 3774 76294
rect 3154 76170 3250 76226
rect 3306 76170 3374 76226
rect 3430 76170 3498 76226
rect 3554 76170 3622 76226
rect 3678 76170 3774 76226
rect 3154 76102 3774 76170
rect 3154 76046 3250 76102
rect 3306 76046 3374 76102
rect 3430 76046 3498 76102
rect 3554 76046 3622 76102
rect 3678 76046 3774 76102
rect 3154 75978 3774 76046
rect 3154 75922 3250 75978
rect 3306 75922 3374 75978
rect 3430 75922 3498 75978
rect 3554 75922 3622 75978
rect 3678 75922 3774 75978
rect 3154 58350 3774 75922
rect 3154 58294 3250 58350
rect 3306 58294 3374 58350
rect 3430 58294 3498 58350
rect 3554 58294 3622 58350
rect 3678 58294 3774 58350
rect 3154 58226 3774 58294
rect 3154 58170 3250 58226
rect 3306 58170 3374 58226
rect 3430 58170 3498 58226
rect 3554 58170 3622 58226
rect 3678 58170 3774 58226
rect 3154 58102 3774 58170
rect 3154 58046 3250 58102
rect 3306 58046 3374 58102
rect 3430 58046 3498 58102
rect 3554 58046 3622 58102
rect 3678 58046 3774 58102
rect 3154 57978 3774 58046
rect 3154 57922 3250 57978
rect 3306 57922 3374 57978
rect 3430 57922 3498 57978
rect 3554 57922 3622 57978
rect 3678 57922 3774 57978
rect 3154 40350 3774 57922
rect 3154 40294 3250 40350
rect 3306 40294 3374 40350
rect 3430 40294 3498 40350
rect 3554 40294 3622 40350
rect 3678 40294 3774 40350
rect 3154 40226 3774 40294
rect 3154 40170 3250 40226
rect 3306 40170 3374 40226
rect 3430 40170 3498 40226
rect 3554 40170 3622 40226
rect 3678 40170 3774 40226
rect 3154 40102 3774 40170
rect 3154 40046 3250 40102
rect 3306 40046 3374 40102
rect 3430 40046 3498 40102
rect 3554 40046 3622 40102
rect 3678 40046 3774 40102
rect 3154 39978 3774 40046
rect 3154 39922 3250 39978
rect 3306 39922 3374 39978
rect 3430 39922 3498 39978
rect 3554 39922 3622 39978
rect 3678 39922 3774 39978
rect 3154 22350 3774 39922
rect 3154 22294 3250 22350
rect 3306 22294 3374 22350
rect 3430 22294 3498 22350
rect 3554 22294 3622 22350
rect 3678 22294 3774 22350
rect 3154 22226 3774 22294
rect 3154 22170 3250 22226
rect 3306 22170 3374 22226
rect 3430 22170 3498 22226
rect 3554 22170 3622 22226
rect 3678 22170 3774 22226
rect 3154 22102 3774 22170
rect 3154 22046 3250 22102
rect 3306 22046 3374 22102
rect 3430 22046 3498 22102
rect 3554 22046 3622 22102
rect 3678 22046 3774 22102
rect 3154 21978 3774 22046
rect 3154 21922 3250 21978
rect 3306 21922 3374 21978
rect 3430 21922 3498 21978
rect 3554 21922 3622 21978
rect 3678 21922 3774 21978
rect 3154 4350 3774 21922
rect 3154 4294 3250 4350
rect 3306 4294 3374 4350
rect 3430 4294 3498 4350
rect 3554 4294 3622 4350
rect 3678 4294 3774 4350
rect 3154 4226 3774 4294
rect 3154 4170 3250 4226
rect 3306 4170 3374 4226
rect 3430 4170 3498 4226
rect 3554 4170 3622 4226
rect 3678 4170 3774 4226
rect 3154 4102 3774 4170
rect 3154 4046 3250 4102
rect 3306 4046 3374 4102
rect 3430 4046 3498 4102
rect 3554 4046 3622 4102
rect 3678 4046 3774 4102
rect 3154 3978 3774 4046
rect 3154 3922 3250 3978
rect 3306 3922 3374 3978
rect 3430 3922 3498 3978
rect 3554 3922 3622 3978
rect 3678 3922 3774 3978
rect 3154 -160 3774 3922
rect 3154 -216 3250 -160
rect 3306 -216 3374 -160
rect 3430 -216 3498 -160
rect 3554 -216 3622 -160
rect 3678 -216 3774 -160
rect 3154 -284 3774 -216
rect 3154 -340 3250 -284
rect 3306 -340 3374 -284
rect 3430 -340 3498 -284
rect 3554 -340 3622 -284
rect 3678 -340 3774 -284
rect 3154 -408 3774 -340
rect 3154 -464 3250 -408
rect 3306 -464 3374 -408
rect 3430 -464 3498 -408
rect 3554 -464 3622 -408
rect 3678 -464 3774 -408
rect 3154 -532 3774 -464
rect 3154 -588 3250 -532
rect 3306 -588 3374 -532
rect 3430 -588 3498 -532
rect 3554 -588 3622 -532
rect 3678 -588 3774 -532
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 -1296 -1120
rect -1916 -1244 -1296 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 -1296 -1244
rect -1916 -1368 -1296 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 -1296 -1368
rect -1916 -1492 -1296 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 -1296 -1492
rect -1916 -1644 -1296 -1548
rect 3154 -1644 3774 -588
rect 6874 598172 7494 598268
rect 6874 598116 6970 598172
rect 7026 598116 7094 598172
rect 7150 598116 7218 598172
rect 7274 598116 7342 598172
rect 7398 598116 7494 598172
rect 6874 598048 7494 598116
rect 6874 597992 6970 598048
rect 7026 597992 7094 598048
rect 7150 597992 7218 598048
rect 7274 597992 7342 598048
rect 7398 597992 7494 598048
rect 6874 597924 7494 597992
rect 6874 597868 6970 597924
rect 7026 597868 7094 597924
rect 7150 597868 7218 597924
rect 7274 597868 7342 597924
rect 7398 597868 7494 597924
rect 6874 597800 7494 597868
rect 6874 597744 6970 597800
rect 7026 597744 7094 597800
rect 7150 597744 7218 597800
rect 7274 597744 7342 597800
rect 7398 597744 7494 597800
rect 6874 586350 7494 597744
rect 6874 586294 6970 586350
rect 7026 586294 7094 586350
rect 7150 586294 7218 586350
rect 7274 586294 7342 586350
rect 7398 586294 7494 586350
rect 6874 586226 7494 586294
rect 6874 586170 6970 586226
rect 7026 586170 7094 586226
rect 7150 586170 7218 586226
rect 7274 586170 7342 586226
rect 7398 586170 7494 586226
rect 6874 586102 7494 586170
rect 6874 586046 6970 586102
rect 7026 586046 7094 586102
rect 7150 586046 7218 586102
rect 7274 586046 7342 586102
rect 7398 586046 7494 586102
rect 6874 585978 7494 586046
rect 6874 585922 6970 585978
rect 7026 585922 7094 585978
rect 7150 585922 7218 585978
rect 7274 585922 7342 585978
rect 7398 585922 7494 585978
rect 6874 568350 7494 585922
rect 6874 568294 6970 568350
rect 7026 568294 7094 568350
rect 7150 568294 7218 568350
rect 7274 568294 7342 568350
rect 7398 568294 7494 568350
rect 6874 568226 7494 568294
rect 6874 568170 6970 568226
rect 7026 568170 7094 568226
rect 7150 568170 7218 568226
rect 7274 568170 7342 568226
rect 7398 568170 7494 568226
rect 6874 568102 7494 568170
rect 6874 568046 6970 568102
rect 7026 568046 7094 568102
rect 7150 568046 7218 568102
rect 7274 568046 7342 568102
rect 7398 568046 7494 568102
rect 6874 567978 7494 568046
rect 6874 567922 6970 567978
rect 7026 567922 7094 567978
rect 7150 567922 7218 567978
rect 7274 567922 7342 567978
rect 7398 567922 7494 567978
rect 6874 550350 7494 567922
rect 6874 550294 6970 550350
rect 7026 550294 7094 550350
rect 7150 550294 7218 550350
rect 7274 550294 7342 550350
rect 7398 550294 7494 550350
rect 6874 550226 7494 550294
rect 6874 550170 6970 550226
rect 7026 550170 7094 550226
rect 7150 550170 7218 550226
rect 7274 550170 7342 550226
rect 7398 550170 7494 550226
rect 6874 550102 7494 550170
rect 6874 550046 6970 550102
rect 7026 550046 7094 550102
rect 7150 550046 7218 550102
rect 7274 550046 7342 550102
rect 7398 550046 7494 550102
rect 6874 549978 7494 550046
rect 6874 549922 6970 549978
rect 7026 549922 7094 549978
rect 7150 549922 7218 549978
rect 7274 549922 7342 549978
rect 7398 549922 7494 549978
rect 6874 532350 7494 549922
rect 6874 532294 6970 532350
rect 7026 532294 7094 532350
rect 7150 532294 7218 532350
rect 7274 532294 7342 532350
rect 7398 532294 7494 532350
rect 6874 532226 7494 532294
rect 6874 532170 6970 532226
rect 7026 532170 7094 532226
rect 7150 532170 7218 532226
rect 7274 532170 7342 532226
rect 7398 532170 7494 532226
rect 6874 532102 7494 532170
rect 6874 532046 6970 532102
rect 7026 532046 7094 532102
rect 7150 532046 7218 532102
rect 7274 532046 7342 532102
rect 7398 532046 7494 532102
rect 6874 531978 7494 532046
rect 6874 531922 6970 531978
rect 7026 531922 7094 531978
rect 7150 531922 7218 531978
rect 7274 531922 7342 531978
rect 7398 531922 7494 531978
rect 6874 514350 7494 531922
rect 6874 514294 6970 514350
rect 7026 514294 7094 514350
rect 7150 514294 7218 514350
rect 7274 514294 7342 514350
rect 7398 514294 7494 514350
rect 6874 514226 7494 514294
rect 6874 514170 6970 514226
rect 7026 514170 7094 514226
rect 7150 514170 7218 514226
rect 7274 514170 7342 514226
rect 7398 514170 7494 514226
rect 6874 514102 7494 514170
rect 6874 514046 6970 514102
rect 7026 514046 7094 514102
rect 7150 514046 7218 514102
rect 7274 514046 7342 514102
rect 7398 514046 7494 514102
rect 6874 513978 7494 514046
rect 6874 513922 6970 513978
rect 7026 513922 7094 513978
rect 7150 513922 7218 513978
rect 7274 513922 7342 513978
rect 7398 513922 7494 513978
rect 6874 496350 7494 513922
rect 6874 496294 6970 496350
rect 7026 496294 7094 496350
rect 7150 496294 7218 496350
rect 7274 496294 7342 496350
rect 7398 496294 7494 496350
rect 6874 496226 7494 496294
rect 6874 496170 6970 496226
rect 7026 496170 7094 496226
rect 7150 496170 7218 496226
rect 7274 496170 7342 496226
rect 7398 496170 7494 496226
rect 6874 496102 7494 496170
rect 6874 496046 6970 496102
rect 7026 496046 7094 496102
rect 7150 496046 7218 496102
rect 7274 496046 7342 496102
rect 7398 496046 7494 496102
rect 6874 495978 7494 496046
rect 6874 495922 6970 495978
rect 7026 495922 7094 495978
rect 7150 495922 7218 495978
rect 7274 495922 7342 495978
rect 7398 495922 7494 495978
rect 6874 478350 7494 495922
rect 6874 478294 6970 478350
rect 7026 478294 7094 478350
rect 7150 478294 7218 478350
rect 7274 478294 7342 478350
rect 7398 478294 7494 478350
rect 6874 478226 7494 478294
rect 6874 478170 6970 478226
rect 7026 478170 7094 478226
rect 7150 478170 7218 478226
rect 7274 478170 7342 478226
rect 7398 478170 7494 478226
rect 6874 478102 7494 478170
rect 6874 478046 6970 478102
rect 7026 478046 7094 478102
rect 7150 478046 7218 478102
rect 7274 478046 7342 478102
rect 7398 478046 7494 478102
rect 6874 477978 7494 478046
rect 6874 477922 6970 477978
rect 7026 477922 7094 477978
rect 7150 477922 7218 477978
rect 7274 477922 7342 477978
rect 7398 477922 7494 477978
rect 6874 460350 7494 477922
rect 6874 460294 6970 460350
rect 7026 460294 7094 460350
rect 7150 460294 7218 460350
rect 7274 460294 7342 460350
rect 7398 460294 7494 460350
rect 6874 460226 7494 460294
rect 6874 460170 6970 460226
rect 7026 460170 7094 460226
rect 7150 460170 7218 460226
rect 7274 460170 7342 460226
rect 7398 460170 7494 460226
rect 6874 460102 7494 460170
rect 6874 460046 6970 460102
rect 7026 460046 7094 460102
rect 7150 460046 7218 460102
rect 7274 460046 7342 460102
rect 7398 460046 7494 460102
rect 6874 459978 7494 460046
rect 6874 459922 6970 459978
rect 7026 459922 7094 459978
rect 7150 459922 7218 459978
rect 7274 459922 7342 459978
rect 7398 459922 7494 459978
rect 6874 442350 7494 459922
rect 6874 442294 6970 442350
rect 7026 442294 7094 442350
rect 7150 442294 7218 442350
rect 7274 442294 7342 442350
rect 7398 442294 7494 442350
rect 6874 442226 7494 442294
rect 6874 442170 6970 442226
rect 7026 442170 7094 442226
rect 7150 442170 7218 442226
rect 7274 442170 7342 442226
rect 7398 442170 7494 442226
rect 6874 442102 7494 442170
rect 6874 442046 6970 442102
rect 7026 442046 7094 442102
rect 7150 442046 7218 442102
rect 7274 442046 7342 442102
rect 7398 442046 7494 442102
rect 6874 441978 7494 442046
rect 6874 441922 6970 441978
rect 7026 441922 7094 441978
rect 7150 441922 7218 441978
rect 7274 441922 7342 441978
rect 7398 441922 7494 441978
rect 6874 424350 7494 441922
rect 6874 424294 6970 424350
rect 7026 424294 7094 424350
rect 7150 424294 7218 424350
rect 7274 424294 7342 424350
rect 7398 424294 7494 424350
rect 6874 424226 7494 424294
rect 6874 424170 6970 424226
rect 7026 424170 7094 424226
rect 7150 424170 7218 424226
rect 7274 424170 7342 424226
rect 7398 424170 7494 424226
rect 6874 424102 7494 424170
rect 6874 424046 6970 424102
rect 7026 424046 7094 424102
rect 7150 424046 7218 424102
rect 7274 424046 7342 424102
rect 7398 424046 7494 424102
rect 6874 423978 7494 424046
rect 6874 423922 6970 423978
rect 7026 423922 7094 423978
rect 7150 423922 7218 423978
rect 7274 423922 7342 423978
rect 7398 423922 7494 423978
rect 6874 406350 7494 423922
rect 6874 406294 6970 406350
rect 7026 406294 7094 406350
rect 7150 406294 7218 406350
rect 7274 406294 7342 406350
rect 7398 406294 7494 406350
rect 6874 406226 7494 406294
rect 6874 406170 6970 406226
rect 7026 406170 7094 406226
rect 7150 406170 7218 406226
rect 7274 406170 7342 406226
rect 7398 406170 7494 406226
rect 6874 406102 7494 406170
rect 6874 406046 6970 406102
rect 7026 406046 7094 406102
rect 7150 406046 7218 406102
rect 7274 406046 7342 406102
rect 7398 406046 7494 406102
rect 6874 405978 7494 406046
rect 6874 405922 6970 405978
rect 7026 405922 7094 405978
rect 7150 405922 7218 405978
rect 7274 405922 7342 405978
rect 7398 405922 7494 405978
rect 6874 388350 7494 405922
rect 6874 388294 6970 388350
rect 7026 388294 7094 388350
rect 7150 388294 7218 388350
rect 7274 388294 7342 388350
rect 7398 388294 7494 388350
rect 6874 388226 7494 388294
rect 6874 388170 6970 388226
rect 7026 388170 7094 388226
rect 7150 388170 7218 388226
rect 7274 388170 7342 388226
rect 7398 388170 7494 388226
rect 6874 388102 7494 388170
rect 6874 388046 6970 388102
rect 7026 388046 7094 388102
rect 7150 388046 7218 388102
rect 7274 388046 7342 388102
rect 7398 388046 7494 388102
rect 6874 387978 7494 388046
rect 6874 387922 6970 387978
rect 7026 387922 7094 387978
rect 7150 387922 7218 387978
rect 7274 387922 7342 387978
rect 7398 387922 7494 387978
rect 6874 370350 7494 387922
rect 6874 370294 6970 370350
rect 7026 370294 7094 370350
rect 7150 370294 7218 370350
rect 7274 370294 7342 370350
rect 7398 370294 7494 370350
rect 6874 370226 7494 370294
rect 6874 370170 6970 370226
rect 7026 370170 7094 370226
rect 7150 370170 7218 370226
rect 7274 370170 7342 370226
rect 7398 370170 7494 370226
rect 6874 370102 7494 370170
rect 6874 370046 6970 370102
rect 7026 370046 7094 370102
rect 7150 370046 7218 370102
rect 7274 370046 7342 370102
rect 7398 370046 7494 370102
rect 6874 369978 7494 370046
rect 6874 369922 6970 369978
rect 7026 369922 7094 369978
rect 7150 369922 7218 369978
rect 7274 369922 7342 369978
rect 7398 369922 7494 369978
rect 6874 352350 7494 369922
rect 6874 352294 6970 352350
rect 7026 352294 7094 352350
rect 7150 352294 7218 352350
rect 7274 352294 7342 352350
rect 7398 352294 7494 352350
rect 6874 352226 7494 352294
rect 6874 352170 6970 352226
rect 7026 352170 7094 352226
rect 7150 352170 7218 352226
rect 7274 352170 7342 352226
rect 7398 352170 7494 352226
rect 6874 352102 7494 352170
rect 6874 352046 6970 352102
rect 7026 352046 7094 352102
rect 7150 352046 7218 352102
rect 7274 352046 7342 352102
rect 7398 352046 7494 352102
rect 6874 351978 7494 352046
rect 6874 351922 6970 351978
rect 7026 351922 7094 351978
rect 7150 351922 7218 351978
rect 7274 351922 7342 351978
rect 7398 351922 7494 351978
rect 6874 334350 7494 351922
rect 6874 334294 6970 334350
rect 7026 334294 7094 334350
rect 7150 334294 7218 334350
rect 7274 334294 7342 334350
rect 7398 334294 7494 334350
rect 6874 334226 7494 334294
rect 6874 334170 6970 334226
rect 7026 334170 7094 334226
rect 7150 334170 7218 334226
rect 7274 334170 7342 334226
rect 7398 334170 7494 334226
rect 6874 334102 7494 334170
rect 6874 334046 6970 334102
rect 7026 334046 7094 334102
rect 7150 334046 7218 334102
rect 7274 334046 7342 334102
rect 7398 334046 7494 334102
rect 6874 333978 7494 334046
rect 6874 333922 6970 333978
rect 7026 333922 7094 333978
rect 7150 333922 7218 333978
rect 7274 333922 7342 333978
rect 7398 333922 7494 333978
rect 6874 316350 7494 333922
rect 6874 316294 6970 316350
rect 7026 316294 7094 316350
rect 7150 316294 7218 316350
rect 7274 316294 7342 316350
rect 7398 316294 7494 316350
rect 6874 316226 7494 316294
rect 6874 316170 6970 316226
rect 7026 316170 7094 316226
rect 7150 316170 7218 316226
rect 7274 316170 7342 316226
rect 7398 316170 7494 316226
rect 6874 316102 7494 316170
rect 6874 316046 6970 316102
rect 7026 316046 7094 316102
rect 7150 316046 7218 316102
rect 7274 316046 7342 316102
rect 7398 316046 7494 316102
rect 6874 315978 7494 316046
rect 6874 315922 6970 315978
rect 7026 315922 7094 315978
rect 7150 315922 7218 315978
rect 7274 315922 7342 315978
rect 7398 315922 7494 315978
rect 6874 298350 7494 315922
rect 6874 298294 6970 298350
rect 7026 298294 7094 298350
rect 7150 298294 7218 298350
rect 7274 298294 7342 298350
rect 7398 298294 7494 298350
rect 6874 298226 7494 298294
rect 6874 298170 6970 298226
rect 7026 298170 7094 298226
rect 7150 298170 7218 298226
rect 7274 298170 7342 298226
rect 7398 298170 7494 298226
rect 6874 298102 7494 298170
rect 6874 298046 6970 298102
rect 7026 298046 7094 298102
rect 7150 298046 7218 298102
rect 7274 298046 7342 298102
rect 7398 298046 7494 298102
rect 6874 297978 7494 298046
rect 6874 297922 6970 297978
rect 7026 297922 7094 297978
rect 7150 297922 7218 297978
rect 7274 297922 7342 297978
rect 7398 297922 7494 297978
rect 6874 280350 7494 297922
rect 6874 280294 6970 280350
rect 7026 280294 7094 280350
rect 7150 280294 7218 280350
rect 7274 280294 7342 280350
rect 7398 280294 7494 280350
rect 6874 280226 7494 280294
rect 6874 280170 6970 280226
rect 7026 280170 7094 280226
rect 7150 280170 7218 280226
rect 7274 280170 7342 280226
rect 7398 280170 7494 280226
rect 6874 280102 7494 280170
rect 6874 280046 6970 280102
rect 7026 280046 7094 280102
rect 7150 280046 7218 280102
rect 7274 280046 7342 280102
rect 7398 280046 7494 280102
rect 6874 279978 7494 280046
rect 6874 279922 6970 279978
rect 7026 279922 7094 279978
rect 7150 279922 7218 279978
rect 7274 279922 7342 279978
rect 7398 279922 7494 279978
rect 6874 262350 7494 279922
rect 6874 262294 6970 262350
rect 7026 262294 7094 262350
rect 7150 262294 7218 262350
rect 7274 262294 7342 262350
rect 7398 262294 7494 262350
rect 6874 262226 7494 262294
rect 6874 262170 6970 262226
rect 7026 262170 7094 262226
rect 7150 262170 7218 262226
rect 7274 262170 7342 262226
rect 7398 262170 7494 262226
rect 6874 262102 7494 262170
rect 6874 262046 6970 262102
rect 7026 262046 7094 262102
rect 7150 262046 7218 262102
rect 7274 262046 7342 262102
rect 7398 262046 7494 262102
rect 6874 261978 7494 262046
rect 6874 261922 6970 261978
rect 7026 261922 7094 261978
rect 7150 261922 7218 261978
rect 7274 261922 7342 261978
rect 7398 261922 7494 261978
rect 6874 244350 7494 261922
rect 6874 244294 6970 244350
rect 7026 244294 7094 244350
rect 7150 244294 7218 244350
rect 7274 244294 7342 244350
rect 7398 244294 7494 244350
rect 6874 244226 7494 244294
rect 6874 244170 6970 244226
rect 7026 244170 7094 244226
rect 7150 244170 7218 244226
rect 7274 244170 7342 244226
rect 7398 244170 7494 244226
rect 6874 244102 7494 244170
rect 6874 244046 6970 244102
rect 7026 244046 7094 244102
rect 7150 244046 7218 244102
rect 7274 244046 7342 244102
rect 7398 244046 7494 244102
rect 6874 243978 7494 244046
rect 6874 243922 6970 243978
rect 7026 243922 7094 243978
rect 7150 243922 7218 243978
rect 7274 243922 7342 243978
rect 7398 243922 7494 243978
rect 6874 226350 7494 243922
rect 6874 226294 6970 226350
rect 7026 226294 7094 226350
rect 7150 226294 7218 226350
rect 7274 226294 7342 226350
rect 7398 226294 7494 226350
rect 6874 226226 7494 226294
rect 6874 226170 6970 226226
rect 7026 226170 7094 226226
rect 7150 226170 7218 226226
rect 7274 226170 7342 226226
rect 7398 226170 7494 226226
rect 6874 226102 7494 226170
rect 6874 226046 6970 226102
rect 7026 226046 7094 226102
rect 7150 226046 7218 226102
rect 7274 226046 7342 226102
rect 7398 226046 7494 226102
rect 6874 225978 7494 226046
rect 6874 225922 6970 225978
rect 7026 225922 7094 225978
rect 7150 225922 7218 225978
rect 7274 225922 7342 225978
rect 7398 225922 7494 225978
rect 6874 208350 7494 225922
rect 6874 208294 6970 208350
rect 7026 208294 7094 208350
rect 7150 208294 7218 208350
rect 7274 208294 7342 208350
rect 7398 208294 7494 208350
rect 6874 208226 7494 208294
rect 6874 208170 6970 208226
rect 7026 208170 7094 208226
rect 7150 208170 7218 208226
rect 7274 208170 7342 208226
rect 7398 208170 7494 208226
rect 6874 208102 7494 208170
rect 6874 208046 6970 208102
rect 7026 208046 7094 208102
rect 7150 208046 7218 208102
rect 7274 208046 7342 208102
rect 7398 208046 7494 208102
rect 6874 207978 7494 208046
rect 6874 207922 6970 207978
rect 7026 207922 7094 207978
rect 7150 207922 7218 207978
rect 7274 207922 7342 207978
rect 7398 207922 7494 207978
rect 6874 190350 7494 207922
rect 6874 190294 6970 190350
rect 7026 190294 7094 190350
rect 7150 190294 7218 190350
rect 7274 190294 7342 190350
rect 7398 190294 7494 190350
rect 6874 190226 7494 190294
rect 6874 190170 6970 190226
rect 7026 190170 7094 190226
rect 7150 190170 7218 190226
rect 7274 190170 7342 190226
rect 7398 190170 7494 190226
rect 6874 190102 7494 190170
rect 6874 190046 6970 190102
rect 7026 190046 7094 190102
rect 7150 190046 7218 190102
rect 7274 190046 7342 190102
rect 7398 190046 7494 190102
rect 6874 189978 7494 190046
rect 6874 189922 6970 189978
rect 7026 189922 7094 189978
rect 7150 189922 7218 189978
rect 7274 189922 7342 189978
rect 7398 189922 7494 189978
rect 6874 172350 7494 189922
rect 6874 172294 6970 172350
rect 7026 172294 7094 172350
rect 7150 172294 7218 172350
rect 7274 172294 7342 172350
rect 7398 172294 7494 172350
rect 6874 172226 7494 172294
rect 6874 172170 6970 172226
rect 7026 172170 7094 172226
rect 7150 172170 7218 172226
rect 7274 172170 7342 172226
rect 7398 172170 7494 172226
rect 6874 172102 7494 172170
rect 6874 172046 6970 172102
rect 7026 172046 7094 172102
rect 7150 172046 7218 172102
rect 7274 172046 7342 172102
rect 7398 172046 7494 172102
rect 6874 171978 7494 172046
rect 6874 171922 6970 171978
rect 7026 171922 7094 171978
rect 7150 171922 7218 171978
rect 7274 171922 7342 171978
rect 7398 171922 7494 171978
rect 6874 154350 7494 171922
rect 6874 154294 6970 154350
rect 7026 154294 7094 154350
rect 7150 154294 7218 154350
rect 7274 154294 7342 154350
rect 7398 154294 7494 154350
rect 6874 154226 7494 154294
rect 6874 154170 6970 154226
rect 7026 154170 7094 154226
rect 7150 154170 7218 154226
rect 7274 154170 7342 154226
rect 7398 154170 7494 154226
rect 6874 154102 7494 154170
rect 6874 154046 6970 154102
rect 7026 154046 7094 154102
rect 7150 154046 7218 154102
rect 7274 154046 7342 154102
rect 7398 154046 7494 154102
rect 6874 153978 7494 154046
rect 6874 153922 6970 153978
rect 7026 153922 7094 153978
rect 7150 153922 7218 153978
rect 7274 153922 7342 153978
rect 7398 153922 7494 153978
rect 6874 136350 7494 153922
rect 6874 136294 6970 136350
rect 7026 136294 7094 136350
rect 7150 136294 7218 136350
rect 7274 136294 7342 136350
rect 7398 136294 7494 136350
rect 6874 136226 7494 136294
rect 6874 136170 6970 136226
rect 7026 136170 7094 136226
rect 7150 136170 7218 136226
rect 7274 136170 7342 136226
rect 7398 136170 7494 136226
rect 6874 136102 7494 136170
rect 6874 136046 6970 136102
rect 7026 136046 7094 136102
rect 7150 136046 7218 136102
rect 7274 136046 7342 136102
rect 7398 136046 7494 136102
rect 6874 135978 7494 136046
rect 6874 135922 6970 135978
rect 7026 135922 7094 135978
rect 7150 135922 7218 135978
rect 7274 135922 7342 135978
rect 7398 135922 7494 135978
rect 6874 118350 7494 135922
rect 6874 118294 6970 118350
rect 7026 118294 7094 118350
rect 7150 118294 7218 118350
rect 7274 118294 7342 118350
rect 7398 118294 7494 118350
rect 6874 118226 7494 118294
rect 6874 118170 6970 118226
rect 7026 118170 7094 118226
rect 7150 118170 7218 118226
rect 7274 118170 7342 118226
rect 7398 118170 7494 118226
rect 6874 118102 7494 118170
rect 6874 118046 6970 118102
rect 7026 118046 7094 118102
rect 7150 118046 7218 118102
rect 7274 118046 7342 118102
rect 7398 118046 7494 118102
rect 6874 117978 7494 118046
rect 6874 117922 6970 117978
rect 7026 117922 7094 117978
rect 7150 117922 7218 117978
rect 7274 117922 7342 117978
rect 7398 117922 7494 117978
rect 6874 100350 7494 117922
rect 6874 100294 6970 100350
rect 7026 100294 7094 100350
rect 7150 100294 7218 100350
rect 7274 100294 7342 100350
rect 7398 100294 7494 100350
rect 6874 100226 7494 100294
rect 6874 100170 6970 100226
rect 7026 100170 7094 100226
rect 7150 100170 7218 100226
rect 7274 100170 7342 100226
rect 7398 100170 7494 100226
rect 6874 100102 7494 100170
rect 6874 100046 6970 100102
rect 7026 100046 7094 100102
rect 7150 100046 7218 100102
rect 7274 100046 7342 100102
rect 7398 100046 7494 100102
rect 6874 99978 7494 100046
rect 6874 99922 6970 99978
rect 7026 99922 7094 99978
rect 7150 99922 7218 99978
rect 7274 99922 7342 99978
rect 7398 99922 7494 99978
rect 6874 82350 7494 99922
rect 6874 82294 6970 82350
rect 7026 82294 7094 82350
rect 7150 82294 7218 82350
rect 7274 82294 7342 82350
rect 7398 82294 7494 82350
rect 6874 82226 7494 82294
rect 6874 82170 6970 82226
rect 7026 82170 7094 82226
rect 7150 82170 7218 82226
rect 7274 82170 7342 82226
rect 7398 82170 7494 82226
rect 6874 82102 7494 82170
rect 6874 82046 6970 82102
rect 7026 82046 7094 82102
rect 7150 82046 7218 82102
rect 7274 82046 7342 82102
rect 7398 82046 7494 82102
rect 6874 81978 7494 82046
rect 6874 81922 6970 81978
rect 7026 81922 7094 81978
rect 7150 81922 7218 81978
rect 7274 81922 7342 81978
rect 7398 81922 7494 81978
rect 6874 64350 7494 81922
rect 6874 64294 6970 64350
rect 7026 64294 7094 64350
rect 7150 64294 7218 64350
rect 7274 64294 7342 64350
rect 7398 64294 7494 64350
rect 6874 64226 7494 64294
rect 6874 64170 6970 64226
rect 7026 64170 7094 64226
rect 7150 64170 7218 64226
rect 7274 64170 7342 64226
rect 7398 64170 7494 64226
rect 6874 64102 7494 64170
rect 6874 64046 6970 64102
rect 7026 64046 7094 64102
rect 7150 64046 7218 64102
rect 7274 64046 7342 64102
rect 7398 64046 7494 64102
rect 6874 63978 7494 64046
rect 6874 63922 6970 63978
rect 7026 63922 7094 63978
rect 7150 63922 7218 63978
rect 7274 63922 7342 63978
rect 7398 63922 7494 63978
rect 6874 46350 7494 63922
rect 6874 46294 6970 46350
rect 7026 46294 7094 46350
rect 7150 46294 7218 46350
rect 7274 46294 7342 46350
rect 7398 46294 7494 46350
rect 6874 46226 7494 46294
rect 6874 46170 6970 46226
rect 7026 46170 7094 46226
rect 7150 46170 7218 46226
rect 7274 46170 7342 46226
rect 7398 46170 7494 46226
rect 6874 46102 7494 46170
rect 6874 46046 6970 46102
rect 7026 46046 7094 46102
rect 7150 46046 7218 46102
rect 7274 46046 7342 46102
rect 7398 46046 7494 46102
rect 6874 45978 7494 46046
rect 6874 45922 6970 45978
rect 7026 45922 7094 45978
rect 7150 45922 7218 45978
rect 7274 45922 7342 45978
rect 7398 45922 7494 45978
rect 6874 28350 7494 45922
rect 6874 28294 6970 28350
rect 7026 28294 7094 28350
rect 7150 28294 7218 28350
rect 7274 28294 7342 28350
rect 7398 28294 7494 28350
rect 6874 28226 7494 28294
rect 6874 28170 6970 28226
rect 7026 28170 7094 28226
rect 7150 28170 7218 28226
rect 7274 28170 7342 28226
rect 7398 28170 7494 28226
rect 6874 28102 7494 28170
rect 6874 28046 6970 28102
rect 7026 28046 7094 28102
rect 7150 28046 7218 28102
rect 7274 28046 7342 28102
rect 7398 28046 7494 28102
rect 6874 27978 7494 28046
rect 6874 27922 6970 27978
rect 7026 27922 7094 27978
rect 7150 27922 7218 27978
rect 7274 27922 7342 27978
rect 7398 27922 7494 27978
rect 6874 10350 7494 27922
rect 6874 10294 6970 10350
rect 7026 10294 7094 10350
rect 7150 10294 7218 10350
rect 7274 10294 7342 10350
rect 7398 10294 7494 10350
rect 6874 10226 7494 10294
rect 6874 10170 6970 10226
rect 7026 10170 7094 10226
rect 7150 10170 7218 10226
rect 7274 10170 7342 10226
rect 7398 10170 7494 10226
rect 6874 10102 7494 10170
rect 6874 10046 6970 10102
rect 7026 10046 7094 10102
rect 7150 10046 7218 10102
rect 7274 10046 7342 10102
rect 7398 10046 7494 10102
rect 6874 9978 7494 10046
rect 6874 9922 6970 9978
rect 7026 9922 7094 9978
rect 7150 9922 7218 9978
rect 7274 9922 7342 9978
rect 7398 9922 7494 9978
rect 6874 -1120 7494 9922
rect 6874 -1176 6970 -1120
rect 7026 -1176 7094 -1120
rect 7150 -1176 7218 -1120
rect 7274 -1176 7342 -1120
rect 7398 -1176 7494 -1120
rect 6874 -1244 7494 -1176
rect 6874 -1300 6970 -1244
rect 7026 -1300 7094 -1244
rect 7150 -1300 7218 -1244
rect 7274 -1300 7342 -1244
rect 7398 -1300 7494 -1244
rect 6874 -1368 7494 -1300
rect 6874 -1424 6970 -1368
rect 7026 -1424 7094 -1368
rect 7150 -1424 7218 -1368
rect 7274 -1424 7342 -1368
rect 7398 -1424 7494 -1368
rect 6874 -1492 7494 -1424
rect 6874 -1548 6970 -1492
rect 7026 -1548 7094 -1492
rect 7150 -1548 7218 -1492
rect 7274 -1548 7342 -1492
rect 7398 -1548 7494 -1492
rect 6874 -1644 7494 -1548
rect 21154 597212 21774 598268
rect 21154 597156 21250 597212
rect 21306 597156 21374 597212
rect 21430 597156 21498 597212
rect 21554 597156 21622 597212
rect 21678 597156 21774 597212
rect 21154 597088 21774 597156
rect 21154 597032 21250 597088
rect 21306 597032 21374 597088
rect 21430 597032 21498 597088
rect 21554 597032 21622 597088
rect 21678 597032 21774 597088
rect 21154 596964 21774 597032
rect 21154 596908 21250 596964
rect 21306 596908 21374 596964
rect 21430 596908 21498 596964
rect 21554 596908 21622 596964
rect 21678 596908 21774 596964
rect 21154 596840 21774 596908
rect 21154 596784 21250 596840
rect 21306 596784 21374 596840
rect 21430 596784 21498 596840
rect 21554 596784 21622 596840
rect 21678 596784 21774 596840
rect 21154 580350 21774 596784
rect 21154 580294 21250 580350
rect 21306 580294 21374 580350
rect 21430 580294 21498 580350
rect 21554 580294 21622 580350
rect 21678 580294 21774 580350
rect 21154 580226 21774 580294
rect 21154 580170 21250 580226
rect 21306 580170 21374 580226
rect 21430 580170 21498 580226
rect 21554 580170 21622 580226
rect 21678 580170 21774 580226
rect 21154 580102 21774 580170
rect 21154 580046 21250 580102
rect 21306 580046 21374 580102
rect 21430 580046 21498 580102
rect 21554 580046 21622 580102
rect 21678 580046 21774 580102
rect 21154 579978 21774 580046
rect 21154 579922 21250 579978
rect 21306 579922 21374 579978
rect 21430 579922 21498 579978
rect 21554 579922 21622 579978
rect 21678 579922 21774 579978
rect 21154 562350 21774 579922
rect 21154 562294 21250 562350
rect 21306 562294 21374 562350
rect 21430 562294 21498 562350
rect 21554 562294 21622 562350
rect 21678 562294 21774 562350
rect 21154 562226 21774 562294
rect 21154 562170 21250 562226
rect 21306 562170 21374 562226
rect 21430 562170 21498 562226
rect 21554 562170 21622 562226
rect 21678 562170 21774 562226
rect 21154 562102 21774 562170
rect 21154 562046 21250 562102
rect 21306 562046 21374 562102
rect 21430 562046 21498 562102
rect 21554 562046 21622 562102
rect 21678 562046 21774 562102
rect 21154 561978 21774 562046
rect 21154 561922 21250 561978
rect 21306 561922 21374 561978
rect 21430 561922 21498 561978
rect 21554 561922 21622 561978
rect 21678 561922 21774 561978
rect 21154 544350 21774 561922
rect 21154 544294 21250 544350
rect 21306 544294 21374 544350
rect 21430 544294 21498 544350
rect 21554 544294 21622 544350
rect 21678 544294 21774 544350
rect 21154 544226 21774 544294
rect 21154 544170 21250 544226
rect 21306 544170 21374 544226
rect 21430 544170 21498 544226
rect 21554 544170 21622 544226
rect 21678 544170 21774 544226
rect 21154 544102 21774 544170
rect 21154 544046 21250 544102
rect 21306 544046 21374 544102
rect 21430 544046 21498 544102
rect 21554 544046 21622 544102
rect 21678 544046 21774 544102
rect 21154 543978 21774 544046
rect 21154 543922 21250 543978
rect 21306 543922 21374 543978
rect 21430 543922 21498 543978
rect 21554 543922 21622 543978
rect 21678 543922 21774 543978
rect 21154 526350 21774 543922
rect 21154 526294 21250 526350
rect 21306 526294 21374 526350
rect 21430 526294 21498 526350
rect 21554 526294 21622 526350
rect 21678 526294 21774 526350
rect 21154 526226 21774 526294
rect 21154 526170 21250 526226
rect 21306 526170 21374 526226
rect 21430 526170 21498 526226
rect 21554 526170 21622 526226
rect 21678 526170 21774 526226
rect 21154 526102 21774 526170
rect 21154 526046 21250 526102
rect 21306 526046 21374 526102
rect 21430 526046 21498 526102
rect 21554 526046 21622 526102
rect 21678 526046 21774 526102
rect 21154 525978 21774 526046
rect 21154 525922 21250 525978
rect 21306 525922 21374 525978
rect 21430 525922 21498 525978
rect 21554 525922 21622 525978
rect 21678 525922 21774 525978
rect 21154 508350 21774 525922
rect 21154 508294 21250 508350
rect 21306 508294 21374 508350
rect 21430 508294 21498 508350
rect 21554 508294 21622 508350
rect 21678 508294 21774 508350
rect 21154 508226 21774 508294
rect 21154 508170 21250 508226
rect 21306 508170 21374 508226
rect 21430 508170 21498 508226
rect 21554 508170 21622 508226
rect 21678 508170 21774 508226
rect 21154 508102 21774 508170
rect 21154 508046 21250 508102
rect 21306 508046 21374 508102
rect 21430 508046 21498 508102
rect 21554 508046 21622 508102
rect 21678 508046 21774 508102
rect 21154 507978 21774 508046
rect 21154 507922 21250 507978
rect 21306 507922 21374 507978
rect 21430 507922 21498 507978
rect 21554 507922 21622 507978
rect 21678 507922 21774 507978
rect 21154 490350 21774 507922
rect 21154 490294 21250 490350
rect 21306 490294 21374 490350
rect 21430 490294 21498 490350
rect 21554 490294 21622 490350
rect 21678 490294 21774 490350
rect 21154 490226 21774 490294
rect 21154 490170 21250 490226
rect 21306 490170 21374 490226
rect 21430 490170 21498 490226
rect 21554 490170 21622 490226
rect 21678 490170 21774 490226
rect 21154 490102 21774 490170
rect 21154 490046 21250 490102
rect 21306 490046 21374 490102
rect 21430 490046 21498 490102
rect 21554 490046 21622 490102
rect 21678 490046 21774 490102
rect 21154 489978 21774 490046
rect 21154 489922 21250 489978
rect 21306 489922 21374 489978
rect 21430 489922 21498 489978
rect 21554 489922 21622 489978
rect 21678 489922 21774 489978
rect 21154 472350 21774 489922
rect 21154 472294 21250 472350
rect 21306 472294 21374 472350
rect 21430 472294 21498 472350
rect 21554 472294 21622 472350
rect 21678 472294 21774 472350
rect 21154 472226 21774 472294
rect 21154 472170 21250 472226
rect 21306 472170 21374 472226
rect 21430 472170 21498 472226
rect 21554 472170 21622 472226
rect 21678 472170 21774 472226
rect 21154 472102 21774 472170
rect 21154 472046 21250 472102
rect 21306 472046 21374 472102
rect 21430 472046 21498 472102
rect 21554 472046 21622 472102
rect 21678 472046 21774 472102
rect 21154 471978 21774 472046
rect 21154 471922 21250 471978
rect 21306 471922 21374 471978
rect 21430 471922 21498 471978
rect 21554 471922 21622 471978
rect 21678 471922 21774 471978
rect 21154 454350 21774 471922
rect 21154 454294 21250 454350
rect 21306 454294 21374 454350
rect 21430 454294 21498 454350
rect 21554 454294 21622 454350
rect 21678 454294 21774 454350
rect 21154 454226 21774 454294
rect 21154 454170 21250 454226
rect 21306 454170 21374 454226
rect 21430 454170 21498 454226
rect 21554 454170 21622 454226
rect 21678 454170 21774 454226
rect 21154 454102 21774 454170
rect 21154 454046 21250 454102
rect 21306 454046 21374 454102
rect 21430 454046 21498 454102
rect 21554 454046 21622 454102
rect 21678 454046 21774 454102
rect 21154 453978 21774 454046
rect 21154 453922 21250 453978
rect 21306 453922 21374 453978
rect 21430 453922 21498 453978
rect 21554 453922 21622 453978
rect 21678 453922 21774 453978
rect 21154 436350 21774 453922
rect 21154 436294 21250 436350
rect 21306 436294 21374 436350
rect 21430 436294 21498 436350
rect 21554 436294 21622 436350
rect 21678 436294 21774 436350
rect 21154 436226 21774 436294
rect 21154 436170 21250 436226
rect 21306 436170 21374 436226
rect 21430 436170 21498 436226
rect 21554 436170 21622 436226
rect 21678 436170 21774 436226
rect 21154 436102 21774 436170
rect 21154 436046 21250 436102
rect 21306 436046 21374 436102
rect 21430 436046 21498 436102
rect 21554 436046 21622 436102
rect 21678 436046 21774 436102
rect 21154 435978 21774 436046
rect 21154 435922 21250 435978
rect 21306 435922 21374 435978
rect 21430 435922 21498 435978
rect 21554 435922 21622 435978
rect 21678 435922 21774 435978
rect 21154 418350 21774 435922
rect 21154 418294 21250 418350
rect 21306 418294 21374 418350
rect 21430 418294 21498 418350
rect 21554 418294 21622 418350
rect 21678 418294 21774 418350
rect 21154 418226 21774 418294
rect 21154 418170 21250 418226
rect 21306 418170 21374 418226
rect 21430 418170 21498 418226
rect 21554 418170 21622 418226
rect 21678 418170 21774 418226
rect 21154 418102 21774 418170
rect 21154 418046 21250 418102
rect 21306 418046 21374 418102
rect 21430 418046 21498 418102
rect 21554 418046 21622 418102
rect 21678 418046 21774 418102
rect 21154 417978 21774 418046
rect 21154 417922 21250 417978
rect 21306 417922 21374 417978
rect 21430 417922 21498 417978
rect 21554 417922 21622 417978
rect 21678 417922 21774 417978
rect 21154 400350 21774 417922
rect 21154 400294 21250 400350
rect 21306 400294 21374 400350
rect 21430 400294 21498 400350
rect 21554 400294 21622 400350
rect 21678 400294 21774 400350
rect 21154 400226 21774 400294
rect 21154 400170 21250 400226
rect 21306 400170 21374 400226
rect 21430 400170 21498 400226
rect 21554 400170 21622 400226
rect 21678 400170 21774 400226
rect 21154 400102 21774 400170
rect 21154 400046 21250 400102
rect 21306 400046 21374 400102
rect 21430 400046 21498 400102
rect 21554 400046 21622 400102
rect 21678 400046 21774 400102
rect 21154 399978 21774 400046
rect 21154 399922 21250 399978
rect 21306 399922 21374 399978
rect 21430 399922 21498 399978
rect 21554 399922 21622 399978
rect 21678 399922 21774 399978
rect 21154 382350 21774 399922
rect 21154 382294 21250 382350
rect 21306 382294 21374 382350
rect 21430 382294 21498 382350
rect 21554 382294 21622 382350
rect 21678 382294 21774 382350
rect 21154 382226 21774 382294
rect 21154 382170 21250 382226
rect 21306 382170 21374 382226
rect 21430 382170 21498 382226
rect 21554 382170 21622 382226
rect 21678 382170 21774 382226
rect 21154 382102 21774 382170
rect 21154 382046 21250 382102
rect 21306 382046 21374 382102
rect 21430 382046 21498 382102
rect 21554 382046 21622 382102
rect 21678 382046 21774 382102
rect 21154 381978 21774 382046
rect 21154 381922 21250 381978
rect 21306 381922 21374 381978
rect 21430 381922 21498 381978
rect 21554 381922 21622 381978
rect 21678 381922 21774 381978
rect 21154 364350 21774 381922
rect 21154 364294 21250 364350
rect 21306 364294 21374 364350
rect 21430 364294 21498 364350
rect 21554 364294 21622 364350
rect 21678 364294 21774 364350
rect 21154 364226 21774 364294
rect 21154 364170 21250 364226
rect 21306 364170 21374 364226
rect 21430 364170 21498 364226
rect 21554 364170 21622 364226
rect 21678 364170 21774 364226
rect 21154 364102 21774 364170
rect 21154 364046 21250 364102
rect 21306 364046 21374 364102
rect 21430 364046 21498 364102
rect 21554 364046 21622 364102
rect 21678 364046 21774 364102
rect 21154 363978 21774 364046
rect 21154 363922 21250 363978
rect 21306 363922 21374 363978
rect 21430 363922 21498 363978
rect 21554 363922 21622 363978
rect 21678 363922 21774 363978
rect 21154 346350 21774 363922
rect 21154 346294 21250 346350
rect 21306 346294 21374 346350
rect 21430 346294 21498 346350
rect 21554 346294 21622 346350
rect 21678 346294 21774 346350
rect 21154 346226 21774 346294
rect 21154 346170 21250 346226
rect 21306 346170 21374 346226
rect 21430 346170 21498 346226
rect 21554 346170 21622 346226
rect 21678 346170 21774 346226
rect 21154 346102 21774 346170
rect 21154 346046 21250 346102
rect 21306 346046 21374 346102
rect 21430 346046 21498 346102
rect 21554 346046 21622 346102
rect 21678 346046 21774 346102
rect 21154 345978 21774 346046
rect 21154 345922 21250 345978
rect 21306 345922 21374 345978
rect 21430 345922 21498 345978
rect 21554 345922 21622 345978
rect 21678 345922 21774 345978
rect 21154 328350 21774 345922
rect 21154 328294 21250 328350
rect 21306 328294 21374 328350
rect 21430 328294 21498 328350
rect 21554 328294 21622 328350
rect 21678 328294 21774 328350
rect 21154 328226 21774 328294
rect 21154 328170 21250 328226
rect 21306 328170 21374 328226
rect 21430 328170 21498 328226
rect 21554 328170 21622 328226
rect 21678 328170 21774 328226
rect 21154 328102 21774 328170
rect 21154 328046 21250 328102
rect 21306 328046 21374 328102
rect 21430 328046 21498 328102
rect 21554 328046 21622 328102
rect 21678 328046 21774 328102
rect 21154 327978 21774 328046
rect 21154 327922 21250 327978
rect 21306 327922 21374 327978
rect 21430 327922 21498 327978
rect 21554 327922 21622 327978
rect 21678 327922 21774 327978
rect 21154 310350 21774 327922
rect 21154 310294 21250 310350
rect 21306 310294 21374 310350
rect 21430 310294 21498 310350
rect 21554 310294 21622 310350
rect 21678 310294 21774 310350
rect 21154 310226 21774 310294
rect 21154 310170 21250 310226
rect 21306 310170 21374 310226
rect 21430 310170 21498 310226
rect 21554 310170 21622 310226
rect 21678 310170 21774 310226
rect 21154 310102 21774 310170
rect 21154 310046 21250 310102
rect 21306 310046 21374 310102
rect 21430 310046 21498 310102
rect 21554 310046 21622 310102
rect 21678 310046 21774 310102
rect 21154 309978 21774 310046
rect 21154 309922 21250 309978
rect 21306 309922 21374 309978
rect 21430 309922 21498 309978
rect 21554 309922 21622 309978
rect 21678 309922 21774 309978
rect 21154 292350 21774 309922
rect 21154 292294 21250 292350
rect 21306 292294 21374 292350
rect 21430 292294 21498 292350
rect 21554 292294 21622 292350
rect 21678 292294 21774 292350
rect 21154 292226 21774 292294
rect 21154 292170 21250 292226
rect 21306 292170 21374 292226
rect 21430 292170 21498 292226
rect 21554 292170 21622 292226
rect 21678 292170 21774 292226
rect 21154 292102 21774 292170
rect 21154 292046 21250 292102
rect 21306 292046 21374 292102
rect 21430 292046 21498 292102
rect 21554 292046 21622 292102
rect 21678 292046 21774 292102
rect 21154 291978 21774 292046
rect 21154 291922 21250 291978
rect 21306 291922 21374 291978
rect 21430 291922 21498 291978
rect 21554 291922 21622 291978
rect 21678 291922 21774 291978
rect 21154 274350 21774 291922
rect 21154 274294 21250 274350
rect 21306 274294 21374 274350
rect 21430 274294 21498 274350
rect 21554 274294 21622 274350
rect 21678 274294 21774 274350
rect 21154 274226 21774 274294
rect 21154 274170 21250 274226
rect 21306 274170 21374 274226
rect 21430 274170 21498 274226
rect 21554 274170 21622 274226
rect 21678 274170 21774 274226
rect 21154 274102 21774 274170
rect 21154 274046 21250 274102
rect 21306 274046 21374 274102
rect 21430 274046 21498 274102
rect 21554 274046 21622 274102
rect 21678 274046 21774 274102
rect 21154 273978 21774 274046
rect 21154 273922 21250 273978
rect 21306 273922 21374 273978
rect 21430 273922 21498 273978
rect 21554 273922 21622 273978
rect 21678 273922 21774 273978
rect 21154 256350 21774 273922
rect 21154 256294 21250 256350
rect 21306 256294 21374 256350
rect 21430 256294 21498 256350
rect 21554 256294 21622 256350
rect 21678 256294 21774 256350
rect 21154 256226 21774 256294
rect 21154 256170 21250 256226
rect 21306 256170 21374 256226
rect 21430 256170 21498 256226
rect 21554 256170 21622 256226
rect 21678 256170 21774 256226
rect 21154 256102 21774 256170
rect 21154 256046 21250 256102
rect 21306 256046 21374 256102
rect 21430 256046 21498 256102
rect 21554 256046 21622 256102
rect 21678 256046 21774 256102
rect 21154 255978 21774 256046
rect 21154 255922 21250 255978
rect 21306 255922 21374 255978
rect 21430 255922 21498 255978
rect 21554 255922 21622 255978
rect 21678 255922 21774 255978
rect 21154 238350 21774 255922
rect 21154 238294 21250 238350
rect 21306 238294 21374 238350
rect 21430 238294 21498 238350
rect 21554 238294 21622 238350
rect 21678 238294 21774 238350
rect 21154 238226 21774 238294
rect 21154 238170 21250 238226
rect 21306 238170 21374 238226
rect 21430 238170 21498 238226
rect 21554 238170 21622 238226
rect 21678 238170 21774 238226
rect 21154 238102 21774 238170
rect 21154 238046 21250 238102
rect 21306 238046 21374 238102
rect 21430 238046 21498 238102
rect 21554 238046 21622 238102
rect 21678 238046 21774 238102
rect 21154 237978 21774 238046
rect 21154 237922 21250 237978
rect 21306 237922 21374 237978
rect 21430 237922 21498 237978
rect 21554 237922 21622 237978
rect 21678 237922 21774 237978
rect 21154 220350 21774 237922
rect 21154 220294 21250 220350
rect 21306 220294 21374 220350
rect 21430 220294 21498 220350
rect 21554 220294 21622 220350
rect 21678 220294 21774 220350
rect 21154 220226 21774 220294
rect 21154 220170 21250 220226
rect 21306 220170 21374 220226
rect 21430 220170 21498 220226
rect 21554 220170 21622 220226
rect 21678 220170 21774 220226
rect 21154 220102 21774 220170
rect 21154 220046 21250 220102
rect 21306 220046 21374 220102
rect 21430 220046 21498 220102
rect 21554 220046 21622 220102
rect 21678 220046 21774 220102
rect 21154 219978 21774 220046
rect 21154 219922 21250 219978
rect 21306 219922 21374 219978
rect 21430 219922 21498 219978
rect 21554 219922 21622 219978
rect 21678 219922 21774 219978
rect 21154 202350 21774 219922
rect 21154 202294 21250 202350
rect 21306 202294 21374 202350
rect 21430 202294 21498 202350
rect 21554 202294 21622 202350
rect 21678 202294 21774 202350
rect 21154 202226 21774 202294
rect 21154 202170 21250 202226
rect 21306 202170 21374 202226
rect 21430 202170 21498 202226
rect 21554 202170 21622 202226
rect 21678 202170 21774 202226
rect 21154 202102 21774 202170
rect 21154 202046 21250 202102
rect 21306 202046 21374 202102
rect 21430 202046 21498 202102
rect 21554 202046 21622 202102
rect 21678 202046 21774 202102
rect 21154 201978 21774 202046
rect 21154 201922 21250 201978
rect 21306 201922 21374 201978
rect 21430 201922 21498 201978
rect 21554 201922 21622 201978
rect 21678 201922 21774 201978
rect 21154 184350 21774 201922
rect 21154 184294 21250 184350
rect 21306 184294 21374 184350
rect 21430 184294 21498 184350
rect 21554 184294 21622 184350
rect 21678 184294 21774 184350
rect 21154 184226 21774 184294
rect 21154 184170 21250 184226
rect 21306 184170 21374 184226
rect 21430 184170 21498 184226
rect 21554 184170 21622 184226
rect 21678 184170 21774 184226
rect 21154 184102 21774 184170
rect 21154 184046 21250 184102
rect 21306 184046 21374 184102
rect 21430 184046 21498 184102
rect 21554 184046 21622 184102
rect 21678 184046 21774 184102
rect 21154 183978 21774 184046
rect 21154 183922 21250 183978
rect 21306 183922 21374 183978
rect 21430 183922 21498 183978
rect 21554 183922 21622 183978
rect 21678 183922 21774 183978
rect 21154 166350 21774 183922
rect 21154 166294 21250 166350
rect 21306 166294 21374 166350
rect 21430 166294 21498 166350
rect 21554 166294 21622 166350
rect 21678 166294 21774 166350
rect 21154 166226 21774 166294
rect 21154 166170 21250 166226
rect 21306 166170 21374 166226
rect 21430 166170 21498 166226
rect 21554 166170 21622 166226
rect 21678 166170 21774 166226
rect 21154 166102 21774 166170
rect 21154 166046 21250 166102
rect 21306 166046 21374 166102
rect 21430 166046 21498 166102
rect 21554 166046 21622 166102
rect 21678 166046 21774 166102
rect 21154 165978 21774 166046
rect 21154 165922 21250 165978
rect 21306 165922 21374 165978
rect 21430 165922 21498 165978
rect 21554 165922 21622 165978
rect 21678 165922 21774 165978
rect 21154 148350 21774 165922
rect 21154 148294 21250 148350
rect 21306 148294 21374 148350
rect 21430 148294 21498 148350
rect 21554 148294 21622 148350
rect 21678 148294 21774 148350
rect 21154 148226 21774 148294
rect 21154 148170 21250 148226
rect 21306 148170 21374 148226
rect 21430 148170 21498 148226
rect 21554 148170 21622 148226
rect 21678 148170 21774 148226
rect 21154 148102 21774 148170
rect 21154 148046 21250 148102
rect 21306 148046 21374 148102
rect 21430 148046 21498 148102
rect 21554 148046 21622 148102
rect 21678 148046 21774 148102
rect 21154 147978 21774 148046
rect 21154 147922 21250 147978
rect 21306 147922 21374 147978
rect 21430 147922 21498 147978
rect 21554 147922 21622 147978
rect 21678 147922 21774 147978
rect 21154 130350 21774 147922
rect 21154 130294 21250 130350
rect 21306 130294 21374 130350
rect 21430 130294 21498 130350
rect 21554 130294 21622 130350
rect 21678 130294 21774 130350
rect 21154 130226 21774 130294
rect 21154 130170 21250 130226
rect 21306 130170 21374 130226
rect 21430 130170 21498 130226
rect 21554 130170 21622 130226
rect 21678 130170 21774 130226
rect 21154 130102 21774 130170
rect 21154 130046 21250 130102
rect 21306 130046 21374 130102
rect 21430 130046 21498 130102
rect 21554 130046 21622 130102
rect 21678 130046 21774 130102
rect 21154 129978 21774 130046
rect 21154 129922 21250 129978
rect 21306 129922 21374 129978
rect 21430 129922 21498 129978
rect 21554 129922 21622 129978
rect 21678 129922 21774 129978
rect 21154 112350 21774 129922
rect 21154 112294 21250 112350
rect 21306 112294 21374 112350
rect 21430 112294 21498 112350
rect 21554 112294 21622 112350
rect 21678 112294 21774 112350
rect 21154 112226 21774 112294
rect 21154 112170 21250 112226
rect 21306 112170 21374 112226
rect 21430 112170 21498 112226
rect 21554 112170 21622 112226
rect 21678 112170 21774 112226
rect 21154 112102 21774 112170
rect 21154 112046 21250 112102
rect 21306 112046 21374 112102
rect 21430 112046 21498 112102
rect 21554 112046 21622 112102
rect 21678 112046 21774 112102
rect 21154 111978 21774 112046
rect 21154 111922 21250 111978
rect 21306 111922 21374 111978
rect 21430 111922 21498 111978
rect 21554 111922 21622 111978
rect 21678 111922 21774 111978
rect 21154 94350 21774 111922
rect 21154 94294 21250 94350
rect 21306 94294 21374 94350
rect 21430 94294 21498 94350
rect 21554 94294 21622 94350
rect 21678 94294 21774 94350
rect 21154 94226 21774 94294
rect 21154 94170 21250 94226
rect 21306 94170 21374 94226
rect 21430 94170 21498 94226
rect 21554 94170 21622 94226
rect 21678 94170 21774 94226
rect 21154 94102 21774 94170
rect 21154 94046 21250 94102
rect 21306 94046 21374 94102
rect 21430 94046 21498 94102
rect 21554 94046 21622 94102
rect 21678 94046 21774 94102
rect 21154 93978 21774 94046
rect 21154 93922 21250 93978
rect 21306 93922 21374 93978
rect 21430 93922 21498 93978
rect 21554 93922 21622 93978
rect 21678 93922 21774 93978
rect 21154 76350 21774 93922
rect 21154 76294 21250 76350
rect 21306 76294 21374 76350
rect 21430 76294 21498 76350
rect 21554 76294 21622 76350
rect 21678 76294 21774 76350
rect 21154 76226 21774 76294
rect 21154 76170 21250 76226
rect 21306 76170 21374 76226
rect 21430 76170 21498 76226
rect 21554 76170 21622 76226
rect 21678 76170 21774 76226
rect 21154 76102 21774 76170
rect 21154 76046 21250 76102
rect 21306 76046 21374 76102
rect 21430 76046 21498 76102
rect 21554 76046 21622 76102
rect 21678 76046 21774 76102
rect 21154 75978 21774 76046
rect 21154 75922 21250 75978
rect 21306 75922 21374 75978
rect 21430 75922 21498 75978
rect 21554 75922 21622 75978
rect 21678 75922 21774 75978
rect 21154 58350 21774 75922
rect 21154 58294 21250 58350
rect 21306 58294 21374 58350
rect 21430 58294 21498 58350
rect 21554 58294 21622 58350
rect 21678 58294 21774 58350
rect 21154 58226 21774 58294
rect 21154 58170 21250 58226
rect 21306 58170 21374 58226
rect 21430 58170 21498 58226
rect 21554 58170 21622 58226
rect 21678 58170 21774 58226
rect 21154 58102 21774 58170
rect 21154 58046 21250 58102
rect 21306 58046 21374 58102
rect 21430 58046 21498 58102
rect 21554 58046 21622 58102
rect 21678 58046 21774 58102
rect 21154 57978 21774 58046
rect 21154 57922 21250 57978
rect 21306 57922 21374 57978
rect 21430 57922 21498 57978
rect 21554 57922 21622 57978
rect 21678 57922 21774 57978
rect 21154 40350 21774 57922
rect 21154 40294 21250 40350
rect 21306 40294 21374 40350
rect 21430 40294 21498 40350
rect 21554 40294 21622 40350
rect 21678 40294 21774 40350
rect 21154 40226 21774 40294
rect 21154 40170 21250 40226
rect 21306 40170 21374 40226
rect 21430 40170 21498 40226
rect 21554 40170 21622 40226
rect 21678 40170 21774 40226
rect 21154 40102 21774 40170
rect 21154 40046 21250 40102
rect 21306 40046 21374 40102
rect 21430 40046 21498 40102
rect 21554 40046 21622 40102
rect 21678 40046 21774 40102
rect 21154 39978 21774 40046
rect 21154 39922 21250 39978
rect 21306 39922 21374 39978
rect 21430 39922 21498 39978
rect 21554 39922 21622 39978
rect 21678 39922 21774 39978
rect 21154 22350 21774 39922
rect 21154 22294 21250 22350
rect 21306 22294 21374 22350
rect 21430 22294 21498 22350
rect 21554 22294 21622 22350
rect 21678 22294 21774 22350
rect 21154 22226 21774 22294
rect 21154 22170 21250 22226
rect 21306 22170 21374 22226
rect 21430 22170 21498 22226
rect 21554 22170 21622 22226
rect 21678 22170 21774 22226
rect 21154 22102 21774 22170
rect 21154 22046 21250 22102
rect 21306 22046 21374 22102
rect 21430 22046 21498 22102
rect 21554 22046 21622 22102
rect 21678 22046 21774 22102
rect 21154 21978 21774 22046
rect 21154 21922 21250 21978
rect 21306 21922 21374 21978
rect 21430 21922 21498 21978
rect 21554 21922 21622 21978
rect 21678 21922 21774 21978
rect 21154 4350 21774 21922
rect 21154 4294 21250 4350
rect 21306 4294 21374 4350
rect 21430 4294 21498 4350
rect 21554 4294 21622 4350
rect 21678 4294 21774 4350
rect 21154 4226 21774 4294
rect 21154 4170 21250 4226
rect 21306 4170 21374 4226
rect 21430 4170 21498 4226
rect 21554 4170 21622 4226
rect 21678 4170 21774 4226
rect 21154 4102 21774 4170
rect 21154 4046 21250 4102
rect 21306 4046 21374 4102
rect 21430 4046 21498 4102
rect 21554 4046 21622 4102
rect 21678 4046 21774 4102
rect 21154 3978 21774 4046
rect 21154 3922 21250 3978
rect 21306 3922 21374 3978
rect 21430 3922 21498 3978
rect 21554 3922 21622 3978
rect 21678 3922 21774 3978
rect 21154 -160 21774 3922
rect 21154 -216 21250 -160
rect 21306 -216 21374 -160
rect 21430 -216 21498 -160
rect 21554 -216 21622 -160
rect 21678 -216 21774 -160
rect 21154 -284 21774 -216
rect 21154 -340 21250 -284
rect 21306 -340 21374 -284
rect 21430 -340 21498 -284
rect 21554 -340 21622 -284
rect 21678 -340 21774 -284
rect 21154 -408 21774 -340
rect 21154 -464 21250 -408
rect 21306 -464 21374 -408
rect 21430 -464 21498 -408
rect 21554 -464 21622 -408
rect 21678 -464 21774 -408
rect 21154 -532 21774 -464
rect 21154 -588 21250 -532
rect 21306 -588 21374 -532
rect 21430 -588 21498 -532
rect 21554 -588 21622 -532
rect 21678 -588 21774 -532
rect 21154 -1644 21774 -588
rect 24874 598172 25494 598268
rect 24874 598116 24970 598172
rect 25026 598116 25094 598172
rect 25150 598116 25218 598172
rect 25274 598116 25342 598172
rect 25398 598116 25494 598172
rect 24874 598048 25494 598116
rect 24874 597992 24970 598048
rect 25026 597992 25094 598048
rect 25150 597992 25218 598048
rect 25274 597992 25342 598048
rect 25398 597992 25494 598048
rect 24874 597924 25494 597992
rect 24874 597868 24970 597924
rect 25026 597868 25094 597924
rect 25150 597868 25218 597924
rect 25274 597868 25342 597924
rect 25398 597868 25494 597924
rect 24874 597800 25494 597868
rect 24874 597744 24970 597800
rect 25026 597744 25094 597800
rect 25150 597744 25218 597800
rect 25274 597744 25342 597800
rect 25398 597744 25494 597800
rect 24874 586350 25494 597744
rect 24874 586294 24970 586350
rect 25026 586294 25094 586350
rect 25150 586294 25218 586350
rect 25274 586294 25342 586350
rect 25398 586294 25494 586350
rect 24874 586226 25494 586294
rect 24874 586170 24970 586226
rect 25026 586170 25094 586226
rect 25150 586170 25218 586226
rect 25274 586170 25342 586226
rect 25398 586170 25494 586226
rect 24874 586102 25494 586170
rect 24874 586046 24970 586102
rect 25026 586046 25094 586102
rect 25150 586046 25218 586102
rect 25274 586046 25342 586102
rect 25398 586046 25494 586102
rect 24874 585978 25494 586046
rect 24874 585922 24970 585978
rect 25026 585922 25094 585978
rect 25150 585922 25218 585978
rect 25274 585922 25342 585978
rect 25398 585922 25494 585978
rect 24874 568350 25494 585922
rect 24874 568294 24970 568350
rect 25026 568294 25094 568350
rect 25150 568294 25218 568350
rect 25274 568294 25342 568350
rect 25398 568294 25494 568350
rect 24874 568226 25494 568294
rect 24874 568170 24970 568226
rect 25026 568170 25094 568226
rect 25150 568170 25218 568226
rect 25274 568170 25342 568226
rect 25398 568170 25494 568226
rect 24874 568102 25494 568170
rect 24874 568046 24970 568102
rect 25026 568046 25094 568102
rect 25150 568046 25218 568102
rect 25274 568046 25342 568102
rect 25398 568046 25494 568102
rect 24874 567978 25494 568046
rect 24874 567922 24970 567978
rect 25026 567922 25094 567978
rect 25150 567922 25218 567978
rect 25274 567922 25342 567978
rect 25398 567922 25494 567978
rect 24874 550350 25494 567922
rect 24874 550294 24970 550350
rect 25026 550294 25094 550350
rect 25150 550294 25218 550350
rect 25274 550294 25342 550350
rect 25398 550294 25494 550350
rect 24874 550226 25494 550294
rect 24874 550170 24970 550226
rect 25026 550170 25094 550226
rect 25150 550170 25218 550226
rect 25274 550170 25342 550226
rect 25398 550170 25494 550226
rect 24874 550102 25494 550170
rect 24874 550046 24970 550102
rect 25026 550046 25094 550102
rect 25150 550046 25218 550102
rect 25274 550046 25342 550102
rect 25398 550046 25494 550102
rect 24874 549978 25494 550046
rect 24874 549922 24970 549978
rect 25026 549922 25094 549978
rect 25150 549922 25218 549978
rect 25274 549922 25342 549978
rect 25398 549922 25494 549978
rect 24874 532350 25494 549922
rect 24874 532294 24970 532350
rect 25026 532294 25094 532350
rect 25150 532294 25218 532350
rect 25274 532294 25342 532350
rect 25398 532294 25494 532350
rect 24874 532226 25494 532294
rect 24874 532170 24970 532226
rect 25026 532170 25094 532226
rect 25150 532170 25218 532226
rect 25274 532170 25342 532226
rect 25398 532170 25494 532226
rect 24874 532102 25494 532170
rect 24874 532046 24970 532102
rect 25026 532046 25094 532102
rect 25150 532046 25218 532102
rect 25274 532046 25342 532102
rect 25398 532046 25494 532102
rect 24874 531978 25494 532046
rect 24874 531922 24970 531978
rect 25026 531922 25094 531978
rect 25150 531922 25218 531978
rect 25274 531922 25342 531978
rect 25398 531922 25494 531978
rect 24874 514350 25494 531922
rect 24874 514294 24970 514350
rect 25026 514294 25094 514350
rect 25150 514294 25218 514350
rect 25274 514294 25342 514350
rect 25398 514294 25494 514350
rect 24874 514226 25494 514294
rect 24874 514170 24970 514226
rect 25026 514170 25094 514226
rect 25150 514170 25218 514226
rect 25274 514170 25342 514226
rect 25398 514170 25494 514226
rect 24874 514102 25494 514170
rect 24874 514046 24970 514102
rect 25026 514046 25094 514102
rect 25150 514046 25218 514102
rect 25274 514046 25342 514102
rect 25398 514046 25494 514102
rect 24874 513978 25494 514046
rect 24874 513922 24970 513978
rect 25026 513922 25094 513978
rect 25150 513922 25218 513978
rect 25274 513922 25342 513978
rect 25398 513922 25494 513978
rect 24874 496350 25494 513922
rect 24874 496294 24970 496350
rect 25026 496294 25094 496350
rect 25150 496294 25218 496350
rect 25274 496294 25342 496350
rect 25398 496294 25494 496350
rect 24874 496226 25494 496294
rect 24874 496170 24970 496226
rect 25026 496170 25094 496226
rect 25150 496170 25218 496226
rect 25274 496170 25342 496226
rect 25398 496170 25494 496226
rect 24874 496102 25494 496170
rect 24874 496046 24970 496102
rect 25026 496046 25094 496102
rect 25150 496046 25218 496102
rect 25274 496046 25342 496102
rect 25398 496046 25494 496102
rect 24874 495978 25494 496046
rect 24874 495922 24970 495978
rect 25026 495922 25094 495978
rect 25150 495922 25218 495978
rect 25274 495922 25342 495978
rect 25398 495922 25494 495978
rect 24874 478350 25494 495922
rect 24874 478294 24970 478350
rect 25026 478294 25094 478350
rect 25150 478294 25218 478350
rect 25274 478294 25342 478350
rect 25398 478294 25494 478350
rect 24874 478226 25494 478294
rect 24874 478170 24970 478226
rect 25026 478170 25094 478226
rect 25150 478170 25218 478226
rect 25274 478170 25342 478226
rect 25398 478170 25494 478226
rect 24874 478102 25494 478170
rect 24874 478046 24970 478102
rect 25026 478046 25094 478102
rect 25150 478046 25218 478102
rect 25274 478046 25342 478102
rect 25398 478046 25494 478102
rect 24874 477978 25494 478046
rect 24874 477922 24970 477978
rect 25026 477922 25094 477978
rect 25150 477922 25218 477978
rect 25274 477922 25342 477978
rect 25398 477922 25494 477978
rect 24874 460350 25494 477922
rect 24874 460294 24970 460350
rect 25026 460294 25094 460350
rect 25150 460294 25218 460350
rect 25274 460294 25342 460350
rect 25398 460294 25494 460350
rect 24874 460226 25494 460294
rect 24874 460170 24970 460226
rect 25026 460170 25094 460226
rect 25150 460170 25218 460226
rect 25274 460170 25342 460226
rect 25398 460170 25494 460226
rect 24874 460102 25494 460170
rect 24874 460046 24970 460102
rect 25026 460046 25094 460102
rect 25150 460046 25218 460102
rect 25274 460046 25342 460102
rect 25398 460046 25494 460102
rect 24874 459978 25494 460046
rect 24874 459922 24970 459978
rect 25026 459922 25094 459978
rect 25150 459922 25218 459978
rect 25274 459922 25342 459978
rect 25398 459922 25494 459978
rect 24874 442350 25494 459922
rect 24874 442294 24970 442350
rect 25026 442294 25094 442350
rect 25150 442294 25218 442350
rect 25274 442294 25342 442350
rect 25398 442294 25494 442350
rect 24874 442226 25494 442294
rect 24874 442170 24970 442226
rect 25026 442170 25094 442226
rect 25150 442170 25218 442226
rect 25274 442170 25342 442226
rect 25398 442170 25494 442226
rect 24874 442102 25494 442170
rect 24874 442046 24970 442102
rect 25026 442046 25094 442102
rect 25150 442046 25218 442102
rect 25274 442046 25342 442102
rect 25398 442046 25494 442102
rect 24874 441978 25494 442046
rect 24874 441922 24970 441978
rect 25026 441922 25094 441978
rect 25150 441922 25218 441978
rect 25274 441922 25342 441978
rect 25398 441922 25494 441978
rect 24874 424350 25494 441922
rect 24874 424294 24970 424350
rect 25026 424294 25094 424350
rect 25150 424294 25218 424350
rect 25274 424294 25342 424350
rect 25398 424294 25494 424350
rect 24874 424226 25494 424294
rect 24874 424170 24970 424226
rect 25026 424170 25094 424226
rect 25150 424170 25218 424226
rect 25274 424170 25342 424226
rect 25398 424170 25494 424226
rect 24874 424102 25494 424170
rect 24874 424046 24970 424102
rect 25026 424046 25094 424102
rect 25150 424046 25218 424102
rect 25274 424046 25342 424102
rect 25398 424046 25494 424102
rect 24874 423978 25494 424046
rect 24874 423922 24970 423978
rect 25026 423922 25094 423978
rect 25150 423922 25218 423978
rect 25274 423922 25342 423978
rect 25398 423922 25494 423978
rect 24874 406350 25494 423922
rect 24874 406294 24970 406350
rect 25026 406294 25094 406350
rect 25150 406294 25218 406350
rect 25274 406294 25342 406350
rect 25398 406294 25494 406350
rect 24874 406226 25494 406294
rect 24874 406170 24970 406226
rect 25026 406170 25094 406226
rect 25150 406170 25218 406226
rect 25274 406170 25342 406226
rect 25398 406170 25494 406226
rect 24874 406102 25494 406170
rect 24874 406046 24970 406102
rect 25026 406046 25094 406102
rect 25150 406046 25218 406102
rect 25274 406046 25342 406102
rect 25398 406046 25494 406102
rect 24874 405978 25494 406046
rect 24874 405922 24970 405978
rect 25026 405922 25094 405978
rect 25150 405922 25218 405978
rect 25274 405922 25342 405978
rect 25398 405922 25494 405978
rect 24874 388350 25494 405922
rect 24874 388294 24970 388350
rect 25026 388294 25094 388350
rect 25150 388294 25218 388350
rect 25274 388294 25342 388350
rect 25398 388294 25494 388350
rect 24874 388226 25494 388294
rect 24874 388170 24970 388226
rect 25026 388170 25094 388226
rect 25150 388170 25218 388226
rect 25274 388170 25342 388226
rect 25398 388170 25494 388226
rect 24874 388102 25494 388170
rect 24874 388046 24970 388102
rect 25026 388046 25094 388102
rect 25150 388046 25218 388102
rect 25274 388046 25342 388102
rect 25398 388046 25494 388102
rect 24874 387978 25494 388046
rect 24874 387922 24970 387978
rect 25026 387922 25094 387978
rect 25150 387922 25218 387978
rect 25274 387922 25342 387978
rect 25398 387922 25494 387978
rect 24874 370350 25494 387922
rect 24874 370294 24970 370350
rect 25026 370294 25094 370350
rect 25150 370294 25218 370350
rect 25274 370294 25342 370350
rect 25398 370294 25494 370350
rect 24874 370226 25494 370294
rect 24874 370170 24970 370226
rect 25026 370170 25094 370226
rect 25150 370170 25218 370226
rect 25274 370170 25342 370226
rect 25398 370170 25494 370226
rect 24874 370102 25494 370170
rect 24874 370046 24970 370102
rect 25026 370046 25094 370102
rect 25150 370046 25218 370102
rect 25274 370046 25342 370102
rect 25398 370046 25494 370102
rect 24874 369978 25494 370046
rect 24874 369922 24970 369978
rect 25026 369922 25094 369978
rect 25150 369922 25218 369978
rect 25274 369922 25342 369978
rect 25398 369922 25494 369978
rect 24874 352350 25494 369922
rect 24874 352294 24970 352350
rect 25026 352294 25094 352350
rect 25150 352294 25218 352350
rect 25274 352294 25342 352350
rect 25398 352294 25494 352350
rect 24874 352226 25494 352294
rect 24874 352170 24970 352226
rect 25026 352170 25094 352226
rect 25150 352170 25218 352226
rect 25274 352170 25342 352226
rect 25398 352170 25494 352226
rect 24874 352102 25494 352170
rect 24874 352046 24970 352102
rect 25026 352046 25094 352102
rect 25150 352046 25218 352102
rect 25274 352046 25342 352102
rect 25398 352046 25494 352102
rect 24874 351978 25494 352046
rect 24874 351922 24970 351978
rect 25026 351922 25094 351978
rect 25150 351922 25218 351978
rect 25274 351922 25342 351978
rect 25398 351922 25494 351978
rect 24874 334350 25494 351922
rect 24874 334294 24970 334350
rect 25026 334294 25094 334350
rect 25150 334294 25218 334350
rect 25274 334294 25342 334350
rect 25398 334294 25494 334350
rect 24874 334226 25494 334294
rect 24874 334170 24970 334226
rect 25026 334170 25094 334226
rect 25150 334170 25218 334226
rect 25274 334170 25342 334226
rect 25398 334170 25494 334226
rect 24874 334102 25494 334170
rect 24874 334046 24970 334102
rect 25026 334046 25094 334102
rect 25150 334046 25218 334102
rect 25274 334046 25342 334102
rect 25398 334046 25494 334102
rect 24874 333978 25494 334046
rect 24874 333922 24970 333978
rect 25026 333922 25094 333978
rect 25150 333922 25218 333978
rect 25274 333922 25342 333978
rect 25398 333922 25494 333978
rect 24874 316350 25494 333922
rect 24874 316294 24970 316350
rect 25026 316294 25094 316350
rect 25150 316294 25218 316350
rect 25274 316294 25342 316350
rect 25398 316294 25494 316350
rect 24874 316226 25494 316294
rect 24874 316170 24970 316226
rect 25026 316170 25094 316226
rect 25150 316170 25218 316226
rect 25274 316170 25342 316226
rect 25398 316170 25494 316226
rect 24874 316102 25494 316170
rect 24874 316046 24970 316102
rect 25026 316046 25094 316102
rect 25150 316046 25218 316102
rect 25274 316046 25342 316102
rect 25398 316046 25494 316102
rect 24874 315978 25494 316046
rect 24874 315922 24970 315978
rect 25026 315922 25094 315978
rect 25150 315922 25218 315978
rect 25274 315922 25342 315978
rect 25398 315922 25494 315978
rect 24874 298350 25494 315922
rect 24874 298294 24970 298350
rect 25026 298294 25094 298350
rect 25150 298294 25218 298350
rect 25274 298294 25342 298350
rect 25398 298294 25494 298350
rect 24874 298226 25494 298294
rect 24874 298170 24970 298226
rect 25026 298170 25094 298226
rect 25150 298170 25218 298226
rect 25274 298170 25342 298226
rect 25398 298170 25494 298226
rect 24874 298102 25494 298170
rect 24874 298046 24970 298102
rect 25026 298046 25094 298102
rect 25150 298046 25218 298102
rect 25274 298046 25342 298102
rect 25398 298046 25494 298102
rect 24874 297978 25494 298046
rect 24874 297922 24970 297978
rect 25026 297922 25094 297978
rect 25150 297922 25218 297978
rect 25274 297922 25342 297978
rect 25398 297922 25494 297978
rect 24874 280350 25494 297922
rect 24874 280294 24970 280350
rect 25026 280294 25094 280350
rect 25150 280294 25218 280350
rect 25274 280294 25342 280350
rect 25398 280294 25494 280350
rect 24874 280226 25494 280294
rect 24874 280170 24970 280226
rect 25026 280170 25094 280226
rect 25150 280170 25218 280226
rect 25274 280170 25342 280226
rect 25398 280170 25494 280226
rect 24874 280102 25494 280170
rect 24874 280046 24970 280102
rect 25026 280046 25094 280102
rect 25150 280046 25218 280102
rect 25274 280046 25342 280102
rect 25398 280046 25494 280102
rect 24874 279978 25494 280046
rect 24874 279922 24970 279978
rect 25026 279922 25094 279978
rect 25150 279922 25218 279978
rect 25274 279922 25342 279978
rect 25398 279922 25494 279978
rect 24874 262350 25494 279922
rect 24874 262294 24970 262350
rect 25026 262294 25094 262350
rect 25150 262294 25218 262350
rect 25274 262294 25342 262350
rect 25398 262294 25494 262350
rect 24874 262226 25494 262294
rect 24874 262170 24970 262226
rect 25026 262170 25094 262226
rect 25150 262170 25218 262226
rect 25274 262170 25342 262226
rect 25398 262170 25494 262226
rect 24874 262102 25494 262170
rect 24874 262046 24970 262102
rect 25026 262046 25094 262102
rect 25150 262046 25218 262102
rect 25274 262046 25342 262102
rect 25398 262046 25494 262102
rect 24874 261978 25494 262046
rect 24874 261922 24970 261978
rect 25026 261922 25094 261978
rect 25150 261922 25218 261978
rect 25274 261922 25342 261978
rect 25398 261922 25494 261978
rect 24874 244350 25494 261922
rect 24874 244294 24970 244350
rect 25026 244294 25094 244350
rect 25150 244294 25218 244350
rect 25274 244294 25342 244350
rect 25398 244294 25494 244350
rect 24874 244226 25494 244294
rect 24874 244170 24970 244226
rect 25026 244170 25094 244226
rect 25150 244170 25218 244226
rect 25274 244170 25342 244226
rect 25398 244170 25494 244226
rect 24874 244102 25494 244170
rect 24874 244046 24970 244102
rect 25026 244046 25094 244102
rect 25150 244046 25218 244102
rect 25274 244046 25342 244102
rect 25398 244046 25494 244102
rect 24874 243978 25494 244046
rect 24874 243922 24970 243978
rect 25026 243922 25094 243978
rect 25150 243922 25218 243978
rect 25274 243922 25342 243978
rect 25398 243922 25494 243978
rect 24874 226350 25494 243922
rect 24874 226294 24970 226350
rect 25026 226294 25094 226350
rect 25150 226294 25218 226350
rect 25274 226294 25342 226350
rect 25398 226294 25494 226350
rect 24874 226226 25494 226294
rect 24874 226170 24970 226226
rect 25026 226170 25094 226226
rect 25150 226170 25218 226226
rect 25274 226170 25342 226226
rect 25398 226170 25494 226226
rect 24874 226102 25494 226170
rect 24874 226046 24970 226102
rect 25026 226046 25094 226102
rect 25150 226046 25218 226102
rect 25274 226046 25342 226102
rect 25398 226046 25494 226102
rect 24874 225978 25494 226046
rect 24874 225922 24970 225978
rect 25026 225922 25094 225978
rect 25150 225922 25218 225978
rect 25274 225922 25342 225978
rect 25398 225922 25494 225978
rect 24874 208350 25494 225922
rect 24874 208294 24970 208350
rect 25026 208294 25094 208350
rect 25150 208294 25218 208350
rect 25274 208294 25342 208350
rect 25398 208294 25494 208350
rect 24874 208226 25494 208294
rect 24874 208170 24970 208226
rect 25026 208170 25094 208226
rect 25150 208170 25218 208226
rect 25274 208170 25342 208226
rect 25398 208170 25494 208226
rect 24874 208102 25494 208170
rect 24874 208046 24970 208102
rect 25026 208046 25094 208102
rect 25150 208046 25218 208102
rect 25274 208046 25342 208102
rect 25398 208046 25494 208102
rect 24874 207978 25494 208046
rect 24874 207922 24970 207978
rect 25026 207922 25094 207978
rect 25150 207922 25218 207978
rect 25274 207922 25342 207978
rect 25398 207922 25494 207978
rect 24874 190350 25494 207922
rect 24874 190294 24970 190350
rect 25026 190294 25094 190350
rect 25150 190294 25218 190350
rect 25274 190294 25342 190350
rect 25398 190294 25494 190350
rect 24874 190226 25494 190294
rect 24874 190170 24970 190226
rect 25026 190170 25094 190226
rect 25150 190170 25218 190226
rect 25274 190170 25342 190226
rect 25398 190170 25494 190226
rect 24874 190102 25494 190170
rect 24874 190046 24970 190102
rect 25026 190046 25094 190102
rect 25150 190046 25218 190102
rect 25274 190046 25342 190102
rect 25398 190046 25494 190102
rect 24874 189978 25494 190046
rect 24874 189922 24970 189978
rect 25026 189922 25094 189978
rect 25150 189922 25218 189978
rect 25274 189922 25342 189978
rect 25398 189922 25494 189978
rect 24874 172350 25494 189922
rect 24874 172294 24970 172350
rect 25026 172294 25094 172350
rect 25150 172294 25218 172350
rect 25274 172294 25342 172350
rect 25398 172294 25494 172350
rect 24874 172226 25494 172294
rect 24874 172170 24970 172226
rect 25026 172170 25094 172226
rect 25150 172170 25218 172226
rect 25274 172170 25342 172226
rect 25398 172170 25494 172226
rect 24874 172102 25494 172170
rect 24874 172046 24970 172102
rect 25026 172046 25094 172102
rect 25150 172046 25218 172102
rect 25274 172046 25342 172102
rect 25398 172046 25494 172102
rect 24874 171978 25494 172046
rect 24874 171922 24970 171978
rect 25026 171922 25094 171978
rect 25150 171922 25218 171978
rect 25274 171922 25342 171978
rect 25398 171922 25494 171978
rect 24874 154350 25494 171922
rect 24874 154294 24970 154350
rect 25026 154294 25094 154350
rect 25150 154294 25218 154350
rect 25274 154294 25342 154350
rect 25398 154294 25494 154350
rect 24874 154226 25494 154294
rect 24874 154170 24970 154226
rect 25026 154170 25094 154226
rect 25150 154170 25218 154226
rect 25274 154170 25342 154226
rect 25398 154170 25494 154226
rect 24874 154102 25494 154170
rect 24874 154046 24970 154102
rect 25026 154046 25094 154102
rect 25150 154046 25218 154102
rect 25274 154046 25342 154102
rect 25398 154046 25494 154102
rect 24874 153978 25494 154046
rect 24874 153922 24970 153978
rect 25026 153922 25094 153978
rect 25150 153922 25218 153978
rect 25274 153922 25342 153978
rect 25398 153922 25494 153978
rect 24874 136350 25494 153922
rect 24874 136294 24970 136350
rect 25026 136294 25094 136350
rect 25150 136294 25218 136350
rect 25274 136294 25342 136350
rect 25398 136294 25494 136350
rect 24874 136226 25494 136294
rect 24874 136170 24970 136226
rect 25026 136170 25094 136226
rect 25150 136170 25218 136226
rect 25274 136170 25342 136226
rect 25398 136170 25494 136226
rect 24874 136102 25494 136170
rect 24874 136046 24970 136102
rect 25026 136046 25094 136102
rect 25150 136046 25218 136102
rect 25274 136046 25342 136102
rect 25398 136046 25494 136102
rect 24874 135978 25494 136046
rect 24874 135922 24970 135978
rect 25026 135922 25094 135978
rect 25150 135922 25218 135978
rect 25274 135922 25342 135978
rect 25398 135922 25494 135978
rect 24874 118350 25494 135922
rect 24874 118294 24970 118350
rect 25026 118294 25094 118350
rect 25150 118294 25218 118350
rect 25274 118294 25342 118350
rect 25398 118294 25494 118350
rect 24874 118226 25494 118294
rect 24874 118170 24970 118226
rect 25026 118170 25094 118226
rect 25150 118170 25218 118226
rect 25274 118170 25342 118226
rect 25398 118170 25494 118226
rect 24874 118102 25494 118170
rect 24874 118046 24970 118102
rect 25026 118046 25094 118102
rect 25150 118046 25218 118102
rect 25274 118046 25342 118102
rect 25398 118046 25494 118102
rect 24874 117978 25494 118046
rect 24874 117922 24970 117978
rect 25026 117922 25094 117978
rect 25150 117922 25218 117978
rect 25274 117922 25342 117978
rect 25398 117922 25494 117978
rect 24874 100350 25494 117922
rect 24874 100294 24970 100350
rect 25026 100294 25094 100350
rect 25150 100294 25218 100350
rect 25274 100294 25342 100350
rect 25398 100294 25494 100350
rect 24874 100226 25494 100294
rect 24874 100170 24970 100226
rect 25026 100170 25094 100226
rect 25150 100170 25218 100226
rect 25274 100170 25342 100226
rect 25398 100170 25494 100226
rect 24874 100102 25494 100170
rect 24874 100046 24970 100102
rect 25026 100046 25094 100102
rect 25150 100046 25218 100102
rect 25274 100046 25342 100102
rect 25398 100046 25494 100102
rect 24874 99978 25494 100046
rect 24874 99922 24970 99978
rect 25026 99922 25094 99978
rect 25150 99922 25218 99978
rect 25274 99922 25342 99978
rect 25398 99922 25494 99978
rect 24874 82350 25494 99922
rect 24874 82294 24970 82350
rect 25026 82294 25094 82350
rect 25150 82294 25218 82350
rect 25274 82294 25342 82350
rect 25398 82294 25494 82350
rect 24874 82226 25494 82294
rect 24874 82170 24970 82226
rect 25026 82170 25094 82226
rect 25150 82170 25218 82226
rect 25274 82170 25342 82226
rect 25398 82170 25494 82226
rect 24874 82102 25494 82170
rect 24874 82046 24970 82102
rect 25026 82046 25094 82102
rect 25150 82046 25218 82102
rect 25274 82046 25342 82102
rect 25398 82046 25494 82102
rect 24874 81978 25494 82046
rect 24874 81922 24970 81978
rect 25026 81922 25094 81978
rect 25150 81922 25218 81978
rect 25274 81922 25342 81978
rect 25398 81922 25494 81978
rect 24874 64350 25494 81922
rect 24874 64294 24970 64350
rect 25026 64294 25094 64350
rect 25150 64294 25218 64350
rect 25274 64294 25342 64350
rect 25398 64294 25494 64350
rect 24874 64226 25494 64294
rect 24874 64170 24970 64226
rect 25026 64170 25094 64226
rect 25150 64170 25218 64226
rect 25274 64170 25342 64226
rect 25398 64170 25494 64226
rect 24874 64102 25494 64170
rect 24874 64046 24970 64102
rect 25026 64046 25094 64102
rect 25150 64046 25218 64102
rect 25274 64046 25342 64102
rect 25398 64046 25494 64102
rect 24874 63978 25494 64046
rect 24874 63922 24970 63978
rect 25026 63922 25094 63978
rect 25150 63922 25218 63978
rect 25274 63922 25342 63978
rect 25398 63922 25494 63978
rect 24874 46350 25494 63922
rect 24874 46294 24970 46350
rect 25026 46294 25094 46350
rect 25150 46294 25218 46350
rect 25274 46294 25342 46350
rect 25398 46294 25494 46350
rect 24874 46226 25494 46294
rect 24874 46170 24970 46226
rect 25026 46170 25094 46226
rect 25150 46170 25218 46226
rect 25274 46170 25342 46226
rect 25398 46170 25494 46226
rect 24874 46102 25494 46170
rect 24874 46046 24970 46102
rect 25026 46046 25094 46102
rect 25150 46046 25218 46102
rect 25274 46046 25342 46102
rect 25398 46046 25494 46102
rect 24874 45978 25494 46046
rect 24874 45922 24970 45978
rect 25026 45922 25094 45978
rect 25150 45922 25218 45978
rect 25274 45922 25342 45978
rect 25398 45922 25494 45978
rect 24874 28350 25494 45922
rect 24874 28294 24970 28350
rect 25026 28294 25094 28350
rect 25150 28294 25218 28350
rect 25274 28294 25342 28350
rect 25398 28294 25494 28350
rect 24874 28226 25494 28294
rect 24874 28170 24970 28226
rect 25026 28170 25094 28226
rect 25150 28170 25218 28226
rect 25274 28170 25342 28226
rect 25398 28170 25494 28226
rect 24874 28102 25494 28170
rect 24874 28046 24970 28102
rect 25026 28046 25094 28102
rect 25150 28046 25218 28102
rect 25274 28046 25342 28102
rect 25398 28046 25494 28102
rect 24874 27978 25494 28046
rect 24874 27922 24970 27978
rect 25026 27922 25094 27978
rect 25150 27922 25218 27978
rect 25274 27922 25342 27978
rect 25398 27922 25494 27978
rect 24874 10350 25494 27922
rect 24874 10294 24970 10350
rect 25026 10294 25094 10350
rect 25150 10294 25218 10350
rect 25274 10294 25342 10350
rect 25398 10294 25494 10350
rect 24874 10226 25494 10294
rect 24874 10170 24970 10226
rect 25026 10170 25094 10226
rect 25150 10170 25218 10226
rect 25274 10170 25342 10226
rect 25398 10170 25494 10226
rect 24874 10102 25494 10170
rect 24874 10046 24970 10102
rect 25026 10046 25094 10102
rect 25150 10046 25218 10102
rect 25274 10046 25342 10102
rect 25398 10046 25494 10102
rect 24874 9978 25494 10046
rect 24874 9922 24970 9978
rect 25026 9922 25094 9978
rect 25150 9922 25218 9978
rect 25274 9922 25342 9978
rect 25398 9922 25494 9978
rect 24874 -1120 25494 9922
rect 24874 -1176 24970 -1120
rect 25026 -1176 25094 -1120
rect 25150 -1176 25218 -1120
rect 25274 -1176 25342 -1120
rect 25398 -1176 25494 -1120
rect 24874 -1244 25494 -1176
rect 24874 -1300 24970 -1244
rect 25026 -1300 25094 -1244
rect 25150 -1300 25218 -1244
rect 25274 -1300 25342 -1244
rect 25398 -1300 25494 -1244
rect 24874 -1368 25494 -1300
rect 24874 -1424 24970 -1368
rect 25026 -1424 25094 -1368
rect 25150 -1424 25218 -1368
rect 25274 -1424 25342 -1368
rect 25398 -1424 25494 -1368
rect 24874 -1492 25494 -1424
rect 24874 -1548 24970 -1492
rect 25026 -1548 25094 -1492
rect 25150 -1548 25218 -1492
rect 25274 -1548 25342 -1492
rect 25398 -1548 25494 -1492
rect 24874 -1644 25494 -1548
rect 39154 597212 39774 598268
rect 39154 597156 39250 597212
rect 39306 597156 39374 597212
rect 39430 597156 39498 597212
rect 39554 597156 39622 597212
rect 39678 597156 39774 597212
rect 39154 597088 39774 597156
rect 39154 597032 39250 597088
rect 39306 597032 39374 597088
rect 39430 597032 39498 597088
rect 39554 597032 39622 597088
rect 39678 597032 39774 597088
rect 39154 596964 39774 597032
rect 39154 596908 39250 596964
rect 39306 596908 39374 596964
rect 39430 596908 39498 596964
rect 39554 596908 39622 596964
rect 39678 596908 39774 596964
rect 39154 596840 39774 596908
rect 39154 596784 39250 596840
rect 39306 596784 39374 596840
rect 39430 596784 39498 596840
rect 39554 596784 39622 596840
rect 39678 596784 39774 596840
rect 39154 580350 39774 596784
rect 39154 580294 39250 580350
rect 39306 580294 39374 580350
rect 39430 580294 39498 580350
rect 39554 580294 39622 580350
rect 39678 580294 39774 580350
rect 39154 580226 39774 580294
rect 39154 580170 39250 580226
rect 39306 580170 39374 580226
rect 39430 580170 39498 580226
rect 39554 580170 39622 580226
rect 39678 580170 39774 580226
rect 39154 580102 39774 580170
rect 39154 580046 39250 580102
rect 39306 580046 39374 580102
rect 39430 580046 39498 580102
rect 39554 580046 39622 580102
rect 39678 580046 39774 580102
rect 39154 579978 39774 580046
rect 39154 579922 39250 579978
rect 39306 579922 39374 579978
rect 39430 579922 39498 579978
rect 39554 579922 39622 579978
rect 39678 579922 39774 579978
rect 39154 562350 39774 579922
rect 39154 562294 39250 562350
rect 39306 562294 39374 562350
rect 39430 562294 39498 562350
rect 39554 562294 39622 562350
rect 39678 562294 39774 562350
rect 39154 562226 39774 562294
rect 39154 562170 39250 562226
rect 39306 562170 39374 562226
rect 39430 562170 39498 562226
rect 39554 562170 39622 562226
rect 39678 562170 39774 562226
rect 39154 562102 39774 562170
rect 39154 562046 39250 562102
rect 39306 562046 39374 562102
rect 39430 562046 39498 562102
rect 39554 562046 39622 562102
rect 39678 562046 39774 562102
rect 39154 561978 39774 562046
rect 39154 561922 39250 561978
rect 39306 561922 39374 561978
rect 39430 561922 39498 561978
rect 39554 561922 39622 561978
rect 39678 561922 39774 561978
rect 39154 544350 39774 561922
rect 39154 544294 39250 544350
rect 39306 544294 39374 544350
rect 39430 544294 39498 544350
rect 39554 544294 39622 544350
rect 39678 544294 39774 544350
rect 39154 544226 39774 544294
rect 39154 544170 39250 544226
rect 39306 544170 39374 544226
rect 39430 544170 39498 544226
rect 39554 544170 39622 544226
rect 39678 544170 39774 544226
rect 39154 544102 39774 544170
rect 39154 544046 39250 544102
rect 39306 544046 39374 544102
rect 39430 544046 39498 544102
rect 39554 544046 39622 544102
rect 39678 544046 39774 544102
rect 39154 543978 39774 544046
rect 39154 543922 39250 543978
rect 39306 543922 39374 543978
rect 39430 543922 39498 543978
rect 39554 543922 39622 543978
rect 39678 543922 39774 543978
rect 39154 526350 39774 543922
rect 39154 526294 39250 526350
rect 39306 526294 39374 526350
rect 39430 526294 39498 526350
rect 39554 526294 39622 526350
rect 39678 526294 39774 526350
rect 39154 526226 39774 526294
rect 39154 526170 39250 526226
rect 39306 526170 39374 526226
rect 39430 526170 39498 526226
rect 39554 526170 39622 526226
rect 39678 526170 39774 526226
rect 39154 526102 39774 526170
rect 39154 526046 39250 526102
rect 39306 526046 39374 526102
rect 39430 526046 39498 526102
rect 39554 526046 39622 526102
rect 39678 526046 39774 526102
rect 39154 525978 39774 526046
rect 39154 525922 39250 525978
rect 39306 525922 39374 525978
rect 39430 525922 39498 525978
rect 39554 525922 39622 525978
rect 39678 525922 39774 525978
rect 39154 508350 39774 525922
rect 39154 508294 39250 508350
rect 39306 508294 39374 508350
rect 39430 508294 39498 508350
rect 39554 508294 39622 508350
rect 39678 508294 39774 508350
rect 39154 508226 39774 508294
rect 39154 508170 39250 508226
rect 39306 508170 39374 508226
rect 39430 508170 39498 508226
rect 39554 508170 39622 508226
rect 39678 508170 39774 508226
rect 39154 508102 39774 508170
rect 39154 508046 39250 508102
rect 39306 508046 39374 508102
rect 39430 508046 39498 508102
rect 39554 508046 39622 508102
rect 39678 508046 39774 508102
rect 39154 507978 39774 508046
rect 39154 507922 39250 507978
rect 39306 507922 39374 507978
rect 39430 507922 39498 507978
rect 39554 507922 39622 507978
rect 39678 507922 39774 507978
rect 39154 490350 39774 507922
rect 39154 490294 39250 490350
rect 39306 490294 39374 490350
rect 39430 490294 39498 490350
rect 39554 490294 39622 490350
rect 39678 490294 39774 490350
rect 39154 490226 39774 490294
rect 39154 490170 39250 490226
rect 39306 490170 39374 490226
rect 39430 490170 39498 490226
rect 39554 490170 39622 490226
rect 39678 490170 39774 490226
rect 39154 490102 39774 490170
rect 39154 490046 39250 490102
rect 39306 490046 39374 490102
rect 39430 490046 39498 490102
rect 39554 490046 39622 490102
rect 39678 490046 39774 490102
rect 39154 489978 39774 490046
rect 39154 489922 39250 489978
rect 39306 489922 39374 489978
rect 39430 489922 39498 489978
rect 39554 489922 39622 489978
rect 39678 489922 39774 489978
rect 39154 472350 39774 489922
rect 39154 472294 39250 472350
rect 39306 472294 39374 472350
rect 39430 472294 39498 472350
rect 39554 472294 39622 472350
rect 39678 472294 39774 472350
rect 39154 472226 39774 472294
rect 39154 472170 39250 472226
rect 39306 472170 39374 472226
rect 39430 472170 39498 472226
rect 39554 472170 39622 472226
rect 39678 472170 39774 472226
rect 39154 472102 39774 472170
rect 39154 472046 39250 472102
rect 39306 472046 39374 472102
rect 39430 472046 39498 472102
rect 39554 472046 39622 472102
rect 39678 472046 39774 472102
rect 39154 471978 39774 472046
rect 39154 471922 39250 471978
rect 39306 471922 39374 471978
rect 39430 471922 39498 471978
rect 39554 471922 39622 471978
rect 39678 471922 39774 471978
rect 39154 454350 39774 471922
rect 39154 454294 39250 454350
rect 39306 454294 39374 454350
rect 39430 454294 39498 454350
rect 39554 454294 39622 454350
rect 39678 454294 39774 454350
rect 39154 454226 39774 454294
rect 39154 454170 39250 454226
rect 39306 454170 39374 454226
rect 39430 454170 39498 454226
rect 39554 454170 39622 454226
rect 39678 454170 39774 454226
rect 39154 454102 39774 454170
rect 39154 454046 39250 454102
rect 39306 454046 39374 454102
rect 39430 454046 39498 454102
rect 39554 454046 39622 454102
rect 39678 454046 39774 454102
rect 39154 453978 39774 454046
rect 39154 453922 39250 453978
rect 39306 453922 39374 453978
rect 39430 453922 39498 453978
rect 39554 453922 39622 453978
rect 39678 453922 39774 453978
rect 39154 436350 39774 453922
rect 39154 436294 39250 436350
rect 39306 436294 39374 436350
rect 39430 436294 39498 436350
rect 39554 436294 39622 436350
rect 39678 436294 39774 436350
rect 39154 436226 39774 436294
rect 39154 436170 39250 436226
rect 39306 436170 39374 436226
rect 39430 436170 39498 436226
rect 39554 436170 39622 436226
rect 39678 436170 39774 436226
rect 39154 436102 39774 436170
rect 39154 436046 39250 436102
rect 39306 436046 39374 436102
rect 39430 436046 39498 436102
rect 39554 436046 39622 436102
rect 39678 436046 39774 436102
rect 39154 435978 39774 436046
rect 39154 435922 39250 435978
rect 39306 435922 39374 435978
rect 39430 435922 39498 435978
rect 39554 435922 39622 435978
rect 39678 435922 39774 435978
rect 39154 418350 39774 435922
rect 39154 418294 39250 418350
rect 39306 418294 39374 418350
rect 39430 418294 39498 418350
rect 39554 418294 39622 418350
rect 39678 418294 39774 418350
rect 39154 418226 39774 418294
rect 39154 418170 39250 418226
rect 39306 418170 39374 418226
rect 39430 418170 39498 418226
rect 39554 418170 39622 418226
rect 39678 418170 39774 418226
rect 39154 418102 39774 418170
rect 39154 418046 39250 418102
rect 39306 418046 39374 418102
rect 39430 418046 39498 418102
rect 39554 418046 39622 418102
rect 39678 418046 39774 418102
rect 39154 417978 39774 418046
rect 39154 417922 39250 417978
rect 39306 417922 39374 417978
rect 39430 417922 39498 417978
rect 39554 417922 39622 417978
rect 39678 417922 39774 417978
rect 39154 400350 39774 417922
rect 39154 400294 39250 400350
rect 39306 400294 39374 400350
rect 39430 400294 39498 400350
rect 39554 400294 39622 400350
rect 39678 400294 39774 400350
rect 39154 400226 39774 400294
rect 39154 400170 39250 400226
rect 39306 400170 39374 400226
rect 39430 400170 39498 400226
rect 39554 400170 39622 400226
rect 39678 400170 39774 400226
rect 39154 400102 39774 400170
rect 39154 400046 39250 400102
rect 39306 400046 39374 400102
rect 39430 400046 39498 400102
rect 39554 400046 39622 400102
rect 39678 400046 39774 400102
rect 39154 399978 39774 400046
rect 39154 399922 39250 399978
rect 39306 399922 39374 399978
rect 39430 399922 39498 399978
rect 39554 399922 39622 399978
rect 39678 399922 39774 399978
rect 39154 382350 39774 399922
rect 39154 382294 39250 382350
rect 39306 382294 39374 382350
rect 39430 382294 39498 382350
rect 39554 382294 39622 382350
rect 39678 382294 39774 382350
rect 39154 382226 39774 382294
rect 39154 382170 39250 382226
rect 39306 382170 39374 382226
rect 39430 382170 39498 382226
rect 39554 382170 39622 382226
rect 39678 382170 39774 382226
rect 39154 382102 39774 382170
rect 39154 382046 39250 382102
rect 39306 382046 39374 382102
rect 39430 382046 39498 382102
rect 39554 382046 39622 382102
rect 39678 382046 39774 382102
rect 39154 381978 39774 382046
rect 39154 381922 39250 381978
rect 39306 381922 39374 381978
rect 39430 381922 39498 381978
rect 39554 381922 39622 381978
rect 39678 381922 39774 381978
rect 39154 364350 39774 381922
rect 39154 364294 39250 364350
rect 39306 364294 39374 364350
rect 39430 364294 39498 364350
rect 39554 364294 39622 364350
rect 39678 364294 39774 364350
rect 39154 364226 39774 364294
rect 39154 364170 39250 364226
rect 39306 364170 39374 364226
rect 39430 364170 39498 364226
rect 39554 364170 39622 364226
rect 39678 364170 39774 364226
rect 39154 364102 39774 364170
rect 39154 364046 39250 364102
rect 39306 364046 39374 364102
rect 39430 364046 39498 364102
rect 39554 364046 39622 364102
rect 39678 364046 39774 364102
rect 39154 363978 39774 364046
rect 39154 363922 39250 363978
rect 39306 363922 39374 363978
rect 39430 363922 39498 363978
rect 39554 363922 39622 363978
rect 39678 363922 39774 363978
rect 39154 346350 39774 363922
rect 39154 346294 39250 346350
rect 39306 346294 39374 346350
rect 39430 346294 39498 346350
rect 39554 346294 39622 346350
rect 39678 346294 39774 346350
rect 39154 346226 39774 346294
rect 39154 346170 39250 346226
rect 39306 346170 39374 346226
rect 39430 346170 39498 346226
rect 39554 346170 39622 346226
rect 39678 346170 39774 346226
rect 39154 346102 39774 346170
rect 39154 346046 39250 346102
rect 39306 346046 39374 346102
rect 39430 346046 39498 346102
rect 39554 346046 39622 346102
rect 39678 346046 39774 346102
rect 39154 345978 39774 346046
rect 39154 345922 39250 345978
rect 39306 345922 39374 345978
rect 39430 345922 39498 345978
rect 39554 345922 39622 345978
rect 39678 345922 39774 345978
rect 39154 328350 39774 345922
rect 39154 328294 39250 328350
rect 39306 328294 39374 328350
rect 39430 328294 39498 328350
rect 39554 328294 39622 328350
rect 39678 328294 39774 328350
rect 39154 328226 39774 328294
rect 39154 328170 39250 328226
rect 39306 328170 39374 328226
rect 39430 328170 39498 328226
rect 39554 328170 39622 328226
rect 39678 328170 39774 328226
rect 39154 328102 39774 328170
rect 39154 328046 39250 328102
rect 39306 328046 39374 328102
rect 39430 328046 39498 328102
rect 39554 328046 39622 328102
rect 39678 328046 39774 328102
rect 39154 327978 39774 328046
rect 39154 327922 39250 327978
rect 39306 327922 39374 327978
rect 39430 327922 39498 327978
rect 39554 327922 39622 327978
rect 39678 327922 39774 327978
rect 39154 310350 39774 327922
rect 39154 310294 39250 310350
rect 39306 310294 39374 310350
rect 39430 310294 39498 310350
rect 39554 310294 39622 310350
rect 39678 310294 39774 310350
rect 39154 310226 39774 310294
rect 39154 310170 39250 310226
rect 39306 310170 39374 310226
rect 39430 310170 39498 310226
rect 39554 310170 39622 310226
rect 39678 310170 39774 310226
rect 39154 310102 39774 310170
rect 39154 310046 39250 310102
rect 39306 310046 39374 310102
rect 39430 310046 39498 310102
rect 39554 310046 39622 310102
rect 39678 310046 39774 310102
rect 39154 309978 39774 310046
rect 39154 309922 39250 309978
rect 39306 309922 39374 309978
rect 39430 309922 39498 309978
rect 39554 309922 39622 309978
rect 39678 309922 39774 309978
rect 39154 292350 39774 309922
rect 39154 292294 39250 292350
rect 39306 292294 39374 292350
rect 39430 292294 39498 292350
rect 39554 292294 39622 292350
rect 39678 292294 39774 292350
rect 39154 292226 39774 292294
rect 39154 292170 39250 292226
rect 39306 292170 39374 292226
rect 39430 292170 39498 292226
rect 39554 292170 39622 292226
rect 39678 292170 39774 292226
rect 39154 292102 39774 292170
rect 39154 292046 39250 292102
rect 39306 292046 39374 292102
rect 39430 292046 39498 292102
rect 39554 292046 39622 292102
rect 39678 292046 39774 292102
rect 39154 291978 39774 292046
rect 39154 291922 39250 291978
rect 39306 291922 39374 291978
rect 39430 291922 39498 291978
rect 39554 291922 39622 291978
rect 39678 291922 39774 291978
rect 39154 274350 39774 291922
rect 39154 274294 39250 274350
rect 39306 274294 39374 274350
rect 39430 274294 39498 274350
rect 39554 274294 39622 274350
rect 39678 274294 39774 274350
rect 39154 274226 39774 274294
rect 39154 274170 39250 274226
rect 39306 274170 39374 274226
rect 39430 274170 39498 274226
rect 39554 274170 39622 274226
rect 39678 274170 39774 274226
rect 39154 274102 39774 274170
rect 39154 274046 39250 274102
rect 39306 274046 39374 274102
rect 39430 274046 39498 274102
rect 39554 274046 39622 274102
rect 39678 274046 39774 274102
rect 39154 273978 39774 274046
rect 39154 273922 39250 273978
rect 39306 273922 39374 273978
rect 39430 273922 39498 273978
rect 39554 273922 39622 273978
rect 39678 273922 39774 273978
rect 39154 256350 39774 273922
rect 39154 256294 39250 256350
rect 39306 256294 39374 256350
rect 39430 256294 39498 256350
rect 39554 256294 39622 256350
rect 39678 256294 39774 256350
rect 39154 256226 39774 256294
rect 39154 256170 39250 256226
rect 39306 256170 39374 256226
rect 39430 256170 39498 256226
rect 39554 256170 39622 256226
rect 39678 256170 39774 256226
rect 39154 256102 39774 256170
rect 39154 256046 39250 256102
rect 39306 256046 39374 256102
rect 39430 256046 39498 256102
rect 39554 256046 39622 256102
rect 39678 256046 39774 256102
rect 39154 255978 39774 256046
rect 39154 255922 39250 255978
rect 39306 255922 39374 255978
rect 39430 255922 39498 255978
rect 39554 255922 39622 255978
rect 39678 255922 39774 255978
rect 39154 238350 39774 255922
rect 39154 238294 39250 238350
rect 39306 238294 39374 238350
rect 39430 238294 39498 238350
rect 39554 238294 39622 238350
rect 39678 238294 39774 238350
rect 39154 238226 39774 238294
rect 39154 238170 39250 238226
rect 39306 238170 39374 238226
rect 39430 238170 39498 238226
rect 39554 238170 39622 238226
rect 39678 238170 39774 238226
rect 39154 238102 39774 238170
rect 39154 238046 39250 238102
rect 39306 238046 39374 238102
rect 39430 238046 39498 238102
rect 39554 238046 39622 238102
rect 39678 238046 39774 238102
rect 39154 237978 39774 238046
rect 39154 237922 39250 237978
rect 39306 237922 39374 237978
rect 39430 237922 39498 237978
rect 39554 237922 39622 237978
rect 39678 237922 39774 237978
rect 39154 220350 39774 237922
rect 39154 220294 39250 220350
rect 39306 220294 39374 220350
rect 39430 220294 39498 220350
rect 39554 220294 39622 220350
rect 39678 220294 39774 220350
rect 39154 220226 39774 220294
rect 39154 220170 39250 220226
rect 39306 220170 39374 220226
rect 39430 220170 39498 220226
rect 39554 220170 39622 220226
rect 39678 220170 39774 220226
rect 39154 220102 39774 220170
rect 39154 220046 39250 220102
rect 39306 220046 39374 220102
rect 39430 220046 39498 220102
rect 39554 220046 39622 220102
rect 39678 220046 39774 220102
rect 39154 219978 39774 220046
rect 39154 219922 39250 219978
rect 39306 219922 39374 219978
rect 39430 219922 39498 219978
rect 39554 219922 39622 219978
rect 39678 219922 39774 219978
rect 39154 202350 39774 219922
rect 39154 202294 39250 202350
rect 39306 202294 39374 202350
rect 39430 202294 39498 202350
rect 39554 202294 39622 202350
rect 39678 202294 39774 202350
rect 39154 202226 39774 202294
rect 39154 202170 39250 202226
rect 39306 202170 39374 202226
rect 39430 202170 39498 202226
rect 39554 202170 39622 202226
rect 39678 202170 39774 202226
rect 39154 202102 39774 202170
rect 39154 202046 39250 202102
rect 39306 202046 39374 202102
rect 39430 202046 39498 202102
rect 39554 202046 39622 202102
rect 39678 202046 39774 202102
rect 39154 201978 39774 202046
rect 39154 201922 39250 201978
rect 39306 201922 39374 201978
rect 39430 201922 39498 201978
rect 39554 201922 39622 201978
rect 39678 201922 39774 201978
rect 39154 184350 39774 201922
rect 39154 184294 39250 184350
rect 39306 184294 39374 184350
rect 39430 184294 39498 184350
rect 39554 184294 39622 184350
rect 39678 184294 39774 184350
rect 39154 184226 39774 184294
rect 39154 184170 39250 184226
rect 39306 184170 39374 184226
rect 39430 184170 39498 184226
rect 39554 184170 39622 184226
rect 39678 184170 39774 184226
rect 39154 184102 39774 184170
rect 39154 184046 39250 184102
rect 39306 184046 39374 184102
rect 39430 184046 39498 184102
rect 39554 184046 39622 184102
rect 39678 184046 39774 184102
rect 39154 183978 39774 184046
rect 39154 183922 39250 183978
rect 39306 183922 39374 183978
rect 39430 183922 39498 183978
rect 39554 183922 39622 183978
rect 39678 183922 39774 183978
rect 39154 166350 39774 183922
rect 39154 166294 39250 166350
rect 39306 166294 39374 166350
rect 39430 166294 39498 166350
rect 39554 166294 39622 166350
rect 39678 166294 39774 166350
rect 39154 166226 39774 166294
rect 39154 166170 39250 166226
rect 39306 166170 39374 166226
rect 39430 166170 39498 166226
rect 39554 166170 39622 166226
rect 39678 166170 39774 166226
rect 39154 166102 39774 166170
rect 39154 166046 39250 166102
rect 39306 166046 39374 166102
rect 39430 166046 39498 166102
rect 39554 166046 39622 166102
rect 39678 166046 39774 166102
rect 39154 165978 39774 166046
rect 39154 165922 39250 165978
rect 39306 165922 39374 165978
rect 39430 165922 39498 165978
rect 39554 165922 39622 165978
rect 39678 165922 39774 165978
rect 39154 148350 39774 165922
rect 39154 148294 39250 148350
rect 39306 148294 39374 148350
rect 39430 148294 39498 148350
rect 39554 148294 39622 148350
rect 39678 148294 39774 148350
rect 39154 148226 39774 148294
rect 39154 148170 39250 148226
rect 39306 148170 39374 148226
rect 39430 148170 39498 148226
rect 39554 148170 39622 148226
rect 39678 148170 39774 148226
rect 39154 148102 39774 148170
rect 39154 148046 39250 148102
rect 39306 148046 39374 148102
rect 39430 148046 39498 148102
rect 39554 148046 39622 148102
rect 39678 148046 39774 148102
rect 39154 147978 39774 148046
rect 39154 147922 39250 147978
rect 39306 147922 39374 147978
rect 39430 147922 39498 147978
rect 39554 147922 39622 147978
rect 39678 147922 39774 147978
rect 39154 130350 39774 147922
rect 39154 130294 39250 130350
rect 39306 130294 39374 130350
rect 39430 130294 39498 130350
rect 39554 130294 39622 130350
rect 39678 130294 39774 130350
rect 39154 130226 39774 130294
rect 39154 130170 39250 130226
rect 39306 130170 39374 130226
rect 39430 130170 39498 130226
rect 39554 130170 39622 130226
rect 39678 130170 39774 130226
rect 39154 130102 39774 130170
rect 39154 130046 39250 130102
rect 39306 130046 39374 130102
rect 39430 130046 39498 130102
rect 39554 130046 39622 130102
rect 39678 130046 39774 130102
rect 39154 129978 39774 130046
rect 39154 129922 39250 129978
rect 39306 129922 39374 129978
rect 39430 129922 39498 129978
rect 39554 129922 39622 129978
rect 39678 129922 39774 129978
rect 39154 112350 39774 129922
rect 39154 112294 39250 112350
rect 39306 112294 39374 112350
rect 39430 112294 39498 112350
rect 39554 112294 39622 112350
rect 39678 112294 39774 112350
rect 39154 112226 39774 112294
rect 39154 112170 39250 112226
rect 39306 112170 39374 112226
rect 39430 112170 39498 112226
rect 39554 112170 39622 112226
rect 39678 112170 39774 112226
rect 39154 112102 39774 112170
rect 39154 112046 39250 112102
rect 39306 112046 39374 112102
rect 39430 112046 39498 112102
rect 39554 112046 39622 112102
rect 39678 112046 39774 112102
rect 39154 111978 39774 112046
rect 39154 111922 39250 111978
rect 39306 111922 39374 111978
rect 39430 111922 39498 111978
rect 39554 111922 39622 111978
rect 39678 111922 39774 111978
rect 39154 94350 39774 111922
rect 39154 94294 39250 94350
rect 39306 94294 39374 94350
rect 39430 94294 39498 94350
rect 39554 94294 39622 94350
rect 39678 94294 39774 94350
rect 39154 94226 39774 94294
rect 39154 94170 39250 94226
rect 39306 94170 39374 94226
rect 39430 94170 39498 94226
rect 39554 94170 39622 94226
rect 39678 94170 39774 94226
rect 39154 94102 39774 94170
rect 39154 94046 39250 94102
rect 39306 94046 39374 94102
rect 39430 94046 39498 94102
rect 39554 94046 39622 94102
rect 39678 94046 39774 94102
rect 39154 93978 39774 94046
rect 39154 93922 39250 93978
rect 39306 93922 39374 93978
rect 39430 93922 39498 93978
rect 39554 93922 39622 93978
rect 39678 93922 39774 93978
rect 39154 76350 39774 93922
rect 39154 76294 39250 76350
rect 39306 76294 39374 76350
rect 39430 76294 39498 76350
rect 39554 76294 39622 76350
rect 39678 76294 39774 76350
rect 39154 76226 39774 76294
rect 39154 76170 39250 76226
rect 39306 76170 39374 76226
rect 39430 76170 39498 76226
rect 39554 76170 39622 76226
rect 39678 76170 39774 76226
rect 39154 76102 39774 76170
rect 39154 76046 39250 76102
rect 39306 76046 39374 76102
rect 39430 76046 39498 76102
rect 39554 76046 39622 76102
rect 39678 76046 39774 76102
rect 39154 75978 39774 76046
rect 39154 75922 39250 75978
rect 39306 75922 39374 75978
rect 39430 75922 39498 75978
rect 39554 75922 39622 75978
rect 39678 75922 39774 75978
rect 39154 58350 39774 75922
rect 39154 58294 39250 58350
rect 39306 58294 39374 58350
rect 39430 58294 39498 58350
rect 39554 58294 39622 58350
rect 39678 58294 39774 58350
rect 39154 58226 39774 58294
rect 39154 58170 39250 58226
rect 39306 58170 39374 58226
rect 39430 58170 39498 58226
rect 39554 58170 39622 58226
rect 39678 58170 39774 58226
rect 39154 58102 39774 58170
rect 39154 58046 39250 58102
rect 39306 58046 39374 58102
rect 39430 58046 39498 58102
rect 39554 58046 39622 58102
rect 39678 58046 39774 58102
rect 39154 57978 39774 58046
rect 39154 57922 39250 57978
rect 39306 57922 39374 57978
rect 39430 57922 39498 57978
rect 39554 57922 39622 57978
rect 39678 57922 39774 57978
rect 39154 40350 39774 57922
rect 39154 40294 39250 40350
rect 39306 40294 39374 40350
rect 39430 40294 39498 40350
rect 39554 40294 39622 40350
rect 39678 40294 39774 40350
rect 39154 40226 39774 40294
rect 39154 40170 39250 40226
rect 39306 40170 39374 40226
rect 39430 40170 39498 40226
rect 39554 40170 39622 40226
rect 39678 40170 39774 40226
rect 39154 40102 39774 40170
rect 39154 40046 39250 40102
rect 39306 40046 39374 40102
rect 39430 40046 39498 40102
rect 39554 40046 39622 40102
rect 39678 40046 39774 40102
rect 39154 39978 39774 40046
rect 39154 39922 39250 39978
rect 39306 39922 39374 39978
rect 39430 39922 39498 39978
rect 39554 39922 39622 39978
rect 39678 39922 39774 39978
rect 39154 22350 39774 39922
rect 39154 22294 39250 22350
rect 39306 22294 39374 22350
rect 39430 22294 39498 22350
rect 39554 22294 39622 22350
rect 39678 22294 39774 22350
rect 39154 22226 39774 22294
rect 39154 22170 39250 22226
rect 39306 22170 39374 22226
rect 39430 22170 39498 22226
rect 39554 22170 39622 22226
rect 39678 22170 39774 22226
rect 39154 22102 39774 22170
rect 39154 22046 39250 22102
rect 39306 22046 39374 22102
rect 39430 22046 39498 22102
rect 39554 22046 39622 22102
rect 39678 22046 39774 22102
rect 39154 21978 39774 22046
rect 39154 21922 39250 21978
rect 39306 21922 39374 21978
rect 39430 21922 39498 21978
rect 39554 21922 39622 21978
rect 39678 21922 39774 21978
rect 39154 4350 39774 21922
rect 39154 4294 39250 4350
rect 39306 4294 39374 4350
rect 39430 4294 39498 4350
rect 39554 4294 39622 4350
rect 39678 4294 39774 4350
rect 39154 4226 39774 4294
rect 39154 4170 39250 4226
rect 39306 4170 39374 4226
rect 39430 4170 39498 4226
rect 39554 4170 39622 4226
rect 39678 4170 39774 4226
rect 39154 4102 39774 4170
rect 39154 4046 39250 4102
rect 39306 4046 39374 4102
rect 39430 4046 39498 4102
rect 39554 4046 39622 4102
rect 39678 4046 39774 4102
rect 39154 3978 39774 4046
rect 39154 3922 39250 3978
rect 39306 3922 39374 3978
rect 39430 3922 39498 3978
rect 39554 3922 39622 3978
rect 39678 3922 39774 3978
rect 39154 -160 39774 3922
rect 39154 -216 39250 -160
rect 39306 -216 39374 -160
rect 39430 -216 39498 -160
rect 39554 -216 39622 -160
rect 39678 -216 39774 -160
rect 39154 -284 39774 -216
rect 39154 -340 39250 -284
rect 39306 -340 39374 -284
rect 39430 -340 39498 -284
rect 39554 -340 39622 -284
rect 39678 -340 39774 -284
rect 39154 -408 39774 -340
rect 39154 -464 39250 -408
rect 39306 -464 39374 -408
rect 39430 -464 39498 -408
rect 39554 -464 39622 -408
rect 39678 -464 39774 -408
rect 39154 -532 39774 -464
rect 39154 -588 39250 -532
rect 39306 -588 39374 -532
rect 39430 -588 39498 -532
rect 39554 -588 39622 -532
rect 39678 -588 39774 -532
rect 39154 -1644 39774 -588
rect 42874 598172 43494 598268
rect 42874 598116 42970 598172
rect 43026 598116 43094 598172
rect 43150 598116 43218 598172
rect 43274 598116 43342 598172
rect 43398 598116 43494 598172
rect 42874 598048 43494 598116
rect 42874 597992 42970 598048
rect 43026 597992 43094 598048
rect 43150 597992 43218 598048
rect 43274 597992 43342 598048
rect 43398 597992 43494 598048
rect 42874 597924 43494 597992
rect 42874 597868 42970 597924
rect 43026 597868 43094 597924
rect 43150 597868 43218 597924
rect 43274 597868 43342 597924
rect 43398 597868 43494 597924
rect 42874 597800 43494 597868
rect 42874 597744 42970 597800
rect 43026 597744 43094 597800
rect 43150 597744 43218 597800
rect 43274 597744 43342 597800
rect 43398 597744 43494 597800
rect 42874 586350 43494 597744
rect 42874 586294 42970 586350
rect 43026 586294 43094 586350
rect 43150 586294 43218 586350
rect 43274 586294 43342 586350
rect 43398 586294 43494 586350
rect 42874 586226 43494 586294
rect 42874 586170 42970 586226
rect 43026 586170 43094 586226
rect 43150 586170 43218 586226
rect 43274 586170 43342 586226
rect 43398 586170 43494 586226
rect 42874 586102 43494 586170
rect 42874 586046 42970 586102
rect 43026 586046 43094 586102
rect 43150 586046 43218 586102
rect 43274 586046 43342 586102
rect 43398 586046 43494 586102
rect 42874 585978 43494 586046
rect 42874 585922 42970 585978
rect 43026 585922 43094 585978
rect 43150 585922 43218 585978
rect 43274 585922 43342 585978
rect 43398 585922 43494 585978
rect 42874 568350 43494 585922
rect 42874 568294 42970 568350
rect 43026 568294 43094 568350
rect 43150 568294 43218 568350
rect 43274 568294 43342 568350
rect 43398 568294 43494 568350
rect 42874 568226 43494 568294
rect 42874 568170 42970 568226
rect 43026 568170 43094 568226
rect 43150 568170 43218 568226
rect 43274 568170 43342 568226
rect 43398 568170 43494 568226
rect 42874 568102 43494 568170
rect 42874 568046 42970 568102
rect 43026 568046 43094 568102
rect 43150 568046 43218 568102
rect 43274 568046 43342 568102
rect 43398 568046 43494 568102
rect 42874 567978 43494 568046
rect 42874 567922 42970 567978
rect 43026 567922 43094 567978
rect 43150 567922 43218 567978
rect 43274 567922 43342 567978
rect 43398 567922 43494 567978
rect 42874 550350 43494 567922
rect 42874 550294 42970 550350
rect 43026 550294 43094 550350
rect 43150 550294 43218 550350
rect 43274 550294 43342 550350
rect 43398 550294 43494 550350
rect 42874 550226 43494 550294
rect 42874 550170 42970 550226
rect 43026 550170 43094 550226
rect 43150 550170 43218 550226
rect 43274 550170 43342 550226
rect 43398 550170 43494 550226
rect 42874 550102 43494 550170
rect 42874 550046 42970 550102
rect 43026 550046 43094 550102
rect 43150 550046 43218 550102
rect 43274 550046 43342 550102
rect 43398 550046 43494 550102
rect 42874 549978 43494 550046
rect 42874 549922 42970 549978
rect 43026 549922 43094 549978
rect 43150 549922 43218 549978
rect 43274 549922 43342 549978
rect 43398 549922 43494 549978
rect 42874 532350 43494 549922
rect 42874 532294 42970 532350
rect 43026 532294 43094 532350
rect 43150 532294 43218 532350
rect 43274 532294 43342 532350
rect 43398 532294 43494 532350
rect 42874 532226 43494 532294
rect 42874 532170 42970 532226
rect 43026 532170 43094 532226
rect 43150 532170 43218 532226
rect 43274 532170 43342 532226
rect 43398 532170 43494 532226
rect 42874 532102 43494 532170
rect 42874 532046 42970 532102
rect 43026 532046 43094 532102
rect 43150 532046 43218 532102
rect 43274 532046 43342 532102
rect 43398 532046 43494 532102
rect 42874 531978 43494 532046
rect 42874 531922 42970 531978
rect 43026 531922 43094 531978
rect 43150 531922 43218 531978
rect 43274 531922 43342 531978
rect 43398 531922 43494 531978
rect 42874 514350 43494 531922
rect 57154 597212 57774 598268
rect 57154 597156 57250 597212
rect 57306 597156 57374 597212
rect 57430 597156 57498 597212
rect 57554 597156 57622 597212
rect 57678 597156 57774 597212
rect 57154 597088 57774 597156
rect 57154 597032 57250 597088
rect 57306 597032 57374 597088
rect 57430 597032 57498 597088
rect 57554 597032 57622 597088
rect 57678 597032 57774 597088
rect 57154 596964 57774 597032
rect 57154 596908 57250 596964
rect 57306 596908 57374 596964
rect 57430 596908 57498 596964
rect 57554 596908 57622 596964
rect 57678 596908 57774 596964
rect 57154 596840 57774 596908
rect 57154 596784 57250 596840
rect 57306 596784 57374 596840
rect 57430 596784 57498 596840
rect 57554 596784 57622 596840
rect 57678 596784 57774 596840
rect 57154 580350 57774 596784
rect 57154 580294 57250 580350
rect 57306 580294 57374 580350
rect 57430 580294 57498 580350
rect 57554 580294 57622 580350
rect 57678 580294 57774 580350
rect 57154 580226 57774 580294
rect 57154 580170 57250 580226
rect 57306 580170 57374 580226
rect 57430 580170 57498 580226
rect 57554 580170 57622 580226
rect 57678 580170 57774 580226
rect 57154 580102 57774 580170
rect 57154 580046 57250 580102
rect 57306 580046 57374 580102
rect 57430 580046 57498 580102
rect 57554 580046 57622 580102
rect 57678 580046 57774 580102
rect 57154 579978 57774 580046
rect 57154 579922 57250 579978
rect 57306 579922 57374 579978
rect 57430 579922 57498 579978
rect 57554 579922 57622 579978
rect 57678 579922 57774 579978
rect 57154 562350 57774 579922
rect 57154 562294 57250 562350
rect 57306 562294 57374 562350
rect 57430 562294 57498 562350
rect 57554 562294 57622 562350
rect 57678 562294 57774 562350
rect 57154 562226 57774 562294
rect 57154 562170 57250 562226
rect 57306 562170 57374 562226
rect 57430 562170 57498 562226
rect 57554 562170 57622 562226
rect 57678 562170 57774 562226
rect 57154 562102 57774 562170
rect 57154 562046 57250 562102
rect 57306 562046 57374 562102
rect 57430 562046 57498 562102
rect 57554 562046 57622 562102
rect 57678 562046 57774 562102
rect 57154 561978 57774 562046
rect 57154 561922 57250 561978
rect 57306 561922 57374 561978
rect 57430 561922 57498 561978
rect 57554 561922 57622 561978
rect 57678 561922 57774 561978
rect 57154 544350 57774 561922
rect 57154 544294 57250 544350
rect 57306 544294 57374 544350
rect 57430 544294 57498 544350
rect 57554 544294 57622 544350
rect 57678 544294 57774 544350
rect 57154 544226 57774 544294
rect 57154 544170 57250 544226
rect 57306 544170 57374 544226
rect 57430 544170 57498 544226
rect 57554 544170 57622 544226
rect 57678 544170 57774 544226
rect 57154 544102 57774 544170
rect 57154 544046 57250 544102
rect 57306 544046 57374 544102
rect 57430 544046 57498 544102
rect 57554 544046 57622 544102
rect 57678 544046 57774 544102
rect 57154 543978 57774 544046
rect 57154 543922 57250 543978
rect 57306 543922 57374 543978
rect 57430 543922 57498 543978
rect 57554 543922 57622 543978
rect 57678 543922 57774 543978
rect 57154 526350 57774 543922
rect 54448 526293 54768 526332
rect 54448 526237 54518 526293
rect 54574 526237 54642 526293
rect 54698 526237 54768 526293
rect 54448 526169 54768 526237
rect 54448 526113 54518 526169
rect 54574 526113 54642 526169
rect 54698 526113 54768 526169
rect 54448 526045 54768 526113
rect 54448 525989 54518 526045
rect 54574 525989 54642 526045
rect 54698 525989 54768 526045
rect 54448 525921 54768 525989
rect 54448 525865 54518 525921
rect 54574 525865 54642 525921
rect 54698 525865 54768 525921
rect 54448 525826 54768 525865
rect 57154 526294 57250 526350
rect 57306 526294 57374 526350
rect 57430 526294 57498 526350
rect 57554 526294 57622 526350
rect 57678 526294 57774 526350
rect 57154 526226 57774 526294
rect 57154 526170 57250 526226
rect 57306 526170 57374 526226
rect 57430 526170 57498 526226
rect 57554 526170 57622 526226
rect 57678 526170 57774 526226
rect 57154 526102 57774 526170
rect 57154 526046 57250 526102
rect 57306 526046 57374 526102
rect 57430 526046 57498 526102
rect 57554 526046 57622 526102
rect 57678 526046 57774 526102
rect 57154 525978 57774 526046
rect 57154 525922 57250 525978
rect 57306 525922 57374 525978
rect 57430 525922 57498 525978
rect 57554 525922 57622 525978
rect 57678 525922 57774 525978
rect 42874 514294 42970 514350
rect 43026 514294 43094 514350
rect 43150 514294 43218 514350
rect 43274 514294 43342 514350
rect 43398 514294 43494 514350
rect 42874 514226 43494 514294
rect 42874 514170 42970 514226
rect 43026 514170 43094 514226
rect 43150 514170 43218 514226
rect 43274 514170 43342 514226
rect 43398 514170 43494 514226
rect 42874 514102 43494 514170
rect 42874 514046 42970 514102
rect 43026 514046 43094 514102
rect 43150 514046 43218 514102
rect 43274 514046 43342 514102
rect 43398 514046 43494 514102
rect 42874 513978 43494 514046
rect 42874 513922 42970 513978
rect 43026 513922 43094 513978
rect 43150 513922 43218 513978
rect 43274 513922 43342 513978
rect 43398 513922 43494 513978
rect 42874 496350 43494 513922
rect 54448 508350 54768 508384
rect 54448 508294 54518 508350
rect 54574 508294 54642 508350
rect 54698 508294 54768 508350
rect 54448 508226 54768 508294
rect 54448 508170 54518 508226
rect 54574 508170 54642 508226
rect 54698 508170 54768 508226
rect 54448 508102 54768 508170
rect 54448 508046 54518 508102
rect 54574 508046 54642 508102
rect 54698 508046 54768 508102
rect 54448 507978 54768 508046
rect 54448 507922 54518 507978
rect 54574 507922 54642 507978
rect 54698 507922 54768 507978
rect 54448 507888 54768 507922
rect 57154 508350 57774 525922
rect 57154 508294 57250 508350
rect 57306 508294 57374 508350
rect 57430 508294 57498 508350
rect 57554 508294 57622 508350
rect 57678 508294 57774 508350
rect 57154 508226 57774 508294
rect 57154 508170 57250 508226
rect 57306 508170 57374 508226
rect 57430 508170 57498 508226
rect 57554 508170 57622 508226
rect 57678 508170 57774 508226
rect 57154 508102 57774 508170
rect 57154 508046 57250 508102
rect 57306 508046 57374 508102
rect 57430 508046 57498 508102
rect 57554 508046 57622 508102
rect 57678 508046 57774 508102
rect 57154 507978 57774 508046
rect 57154 507922 57250 507978
rect 57306 507922 57374 507978
rect 57430 507922 57498 507978
rect 57554 507922 57622 507978
rect 57678 507922 57774 507978
rect 42874 496294 42970 496350
rect 43026 496294 43094 496350
rect 43150 496294 43218 496350
rect 43274 496294 43342 496350
rect 43398 496294 43494 496350
rect 42874 496226 43494 496294
rect 42874 496170 42970 496226
rect 43026 496170 43094 496226
rect 43150 496170 43218 496226
rect 43274 496170 43342 496226
rect 43398 496170 43494 496226
rect 42874 496102 43494 496170
rect 42874 496046 42970 496102
rect 43026 496046 43094 496102
rect 43150 496046 43218 496102
rect 43274 496046 43342 496102
rect 43398 496046 43494 496102
rect 42874 495978 43494 496046
rect 42874 495922 42970 495978
rect 43026 495922 43094 495978
rect 43150 495922 43218 495978
rect 43274 495922 43342 495978
rect 43398 495922 43494 495978
rect 42874 478350 43494 495922
rect 54448 490350 54768 490384
rect 54448 490294 54518 490350
rect 54574 490294 54642 490350
rect 54698 490294 54768 490350
rect 54448 490226 54768 490294
rect 54448 490170 54518 490226
rect 54574 490170 54642 490226
rect 54698 490170 54768 490226
rect 54448 490102 54768 490170
rect 54448 490046 54518 490102
rect 54574 490046 54642 490102
rect 54698 490046 54768 490102
rect 54448 489978 54768 490046
rect 54448 489922 54518 489978
rect 54574 489922 54642 489978
rect 54698 489922 54768 489978
rect 54448 489888 54768 489922
rect 57154 490350 57774 507922
rect 57154 490294 57250 490350
rect 57306 490294 57374 490350
rect 57430 490294 57498 490350
rect 57554 490294 57622 490350
rect 57678 490294 57774 490350
rect 57154 490226 57774 490294
rect 57154 490170 57250 490226
rect 57306 490170 57374 490226
rect 57430 490170 57498 490226
rect 57554 490170 57622 490226
rect 57678 490170 57774 490226
rect 57154 490102 57774 490170
rect 57154 490046 57250 490102
rect 57306 490046 57374 490102
rect 57430 490046 57498 490102
rect 57554 490046 57622 490102
rect 57678 490046 57774 490102
rect 57154 489978 57774 490046
rect 57154 489922 57250 489978
rect 57306 489922 57374 489978
rect 57430 489922 57498 489978
rect 57554 489922 57622 489978
rect 57678 489922 57774 489978
rect 42874 478294 42970 478350
rect 43026 478294 43094 478350
rect 43150 478294 43218 478350
rect 43274 478294 43342 478350
rect 43398 478294 43494 478350
rect 42874 478226 43494 478294
rect 42874 478170 42970 478226
rect 43026 478170 43094 478226
rect 43150 478170 43218 478226
rect 43274 478170 43342 478226
rect 43398 478170 43494 478226
rect 42874 478102 43494 478170
rect 42874 478046 42970 478102
rect 43026 478046 43094 478102
rect 43150 478046 43218 478102
rect 43274 478046 43342 478102
rect 43398 478046 43494 478102
rect 42874 477978 43494 478046
rect 42874 477922 42970 477978
rect 43026 477922 43094 477978
rect 43150 477922 43218 477978
rect 43274 477922 43342 477978
rect 43398 477922 43494 477978
rect 42874 460350 43494 477922
rect 54448 472350 54768 472384
rect 54448 472294 54518 472350
rect 54574 472294 54642 472350
rect 54698 472294 54768 472350
rect 54448 472226 54768 472294
rect 54448 472170 54518 472226
rect 54574 472170 54642 472226
rect 54698 472170 54768 472226
rect 54448 472102 54768 472170
rect 54448 472046 54518 472102
rect 54574 472046 54642 472102
rect 54698 472046 54768 472102
rect 54448 471978 54768 472046
rect 54448 471922 54518 471978
rect 54574 471922 54642 471978
rect 54698 471922 54768 471978
rect 54448 471888 54768 471922
rect 57154 472350 57774 489922
rect 57154 472294 57250 472350
rect 57306 472294 57374 472350
rect 57430 472294 57498 472350
rect 57554 472294 57622 472350
rect 57678 472294 57774 472350
rect 57154 472226 57774 472294
rect 57154 472170 57250 472226
rect 57306 472170 57374 472226
rect 57430 472170 57498 472226
rect 57554 472170 57622 472226
rect 57678 472170 57774 472226
rect 57154 472102 57774 472170
rect 57154 472046 57250 472102
rect 57306 472046 57374 472102
rect 57430 472046 57498 472102
rect 57554 472046 57622 472102
rect 57678 472046 57774 472102
rect 57154 471978 57774 472046
rect 57154 471922 57250 471978
rect 57306 471922 57374 471978
rect 57430 471922 57498 471978
rect 57554 471922 57622 471978
rect 57678 471922 57774 471978
rect 42874 460294 42970 460350
rect 43026 460294 43094 460350
rect 43150 460294 43218 460350
rect 43274 460294 43342 460350
rect 43398 460294 43494 460350
rect 42874 460226 43494 460294
rect 42874 460170 42970 460226
rect 43026 460170 43094 460226
rect 43150 460170 43218 460226
rect 43274 460170 43342 460226
rect 43398 460170 43494 460226
rect 42874 460102 43494 460170
rect 42874 460046 42970 460102
rect 43026 460046 43094 460102
rect 43150 460046 43218 460102
rect 43274 460046 43342 460102
rect 43398 460046 43494 460102
rect 42874 459978 43494 460046
rect 42874 459922 42970 459978
rect 43026 459922 43094 459978
rect 43150 459922 43218 459978
rect 43274 459922 43342 459978
rect 43398 459922 43494 459978
rect 42874 442350 43494 459922
rect 54448 454350 54768 454384
rect 54448 454294 54518 454350
rect 54574 454294 54642 454350
rect 54698 454294 54768 454350
rect 54448 454226 54768 454294
rect 54448 454170 54518 454226
rect 54574 454170 54642 454226
rect 54698 454170 54768 454226
rect 54448 454102 54768 454170
rect 54448 454046 54518 454102
rect 54574 454046 54642 454102
rect 54698 454046 54768 454102
rect 54448 453978 54768 454046
rect 54448 453922 54518 453978
rect 54574 453922 54642 453978
rect 54698 453922 54768 453978
rect 54448 453888 54768 453922
rect 57154 454350 57774 471922
rect 57154 454294 57250 454350
rect 57306 454294 57374 454350
rect 57430 454294 57498 454350
rect 57554 454294 57622 454350
rect 57678 454294 57774 454350
rect 57154 454226 57774 454294
rect 57154 454170 57250 454226
rect 57306 454170 57374 454226
rect 57430 454170 57498 454226
rect 57554 454170 57622 454226
rect 57678 454170 57774 454226
rect 57154 454102 57774 454170
rect 57154 454046 57250 454102
rect 57306 454046 57374 454102
rect 57430 454046 57498 454102
rect 57554 454046 57622 454102
rect 57678 454046 57774 454102
rect 57154 453978 57774 454046
rect 57154 453922 57250 453978
rect 57306 453922 57374 453978
rect 57430 453922 57498 453978
rect 57554 453922 57622 453978
rect 57678 453922 57774 453978
rect 42874 442294 42970 442350
rect 43026 442294 43094 442350
rect 43150 442294 43218 442350
rect 43274 442294 43342 442350
rect 43398 442294 43494 442350
rect 42874 442226 43494 442294
rect 42874 442170 42970 442226
rect 43026 442170 43094 442226
rect 43150 442170 43218 442226
rect 43274 442170 43342 442226
rect 43398 442170 43494 442226
rect 42874 442102 43494 442170
rect 42874 442046 42970 442102
rect 43026 442046 43094 442102
rect 43150 442046 43218 442102
rect 43274 442046 43342 442102
rect 43398 442046 43494 442102
rect 42874 441978 43494 442046
rect 42874 441922 42970 441978
rect 43026 441922 43094 441978
rect 43150 441922 43218 441978
rect 43274 441922 43342 441978
rect 43398 441922 43494 441978
rect 42874 424350 43494 441922
rect 54448 436350 54768 436384
rect 54448 436294 54518 436350
rect 54574 436294 54642 436350
rect 54698 436294 54768 436350
rect 54448 436226 54768 436294
rect 54448 436170 54518 436226
rect 54574 436170 54642 436226
rect 54698 436170 54768 436226
rect 54448 436102 54768 436170
rect 54448 436046 54518 436102
rect 54574 436046 54642 436102
rect 54698 436046 54768 436102
rect 54448 435978 54768 436046
rect 54448 435922 54518 435978
rect 54574 435922 54642 435978
rect 54698 435922 54768 435978
rect 54448 435888 54768 435922
rect 57154 436350 57774 453922
rect 57154 436294 57250 436350
rect 57306 436294 57374 436350
rect 57430 436294 57498 436350
rect 57554 436294 57622 436350
rect 57678 436294 57774 436350
rect 57154 436226 57774 436294
rect 57154 436170 57250 436226
rect 57306 436170 57374 436226
rect 57430 436170 57498 436226
rect 57554 436170 57622 436226
rect 57678 436170 57774 436226
rect 57154 436102 57774 436170
rect 57154 436046 57250 436102
rect 57306 436046 57374 436102
rect 57430 436046 57498 436102
rect 57554 436046 57622 436102
rect 57678 436046 57774 436102
rect 57154 435978 57774 436046
rect 57154 435922 57250 435978
rect 57306 435922 57374 435978
rect 57430 435922 57498 435978
rect 57554 435922 57622 435978
rect 57678 435922 57774 435978
rect 42874 424294 42970 424350
rect 43026 424294 43094 424350
rect 43150 424294 43218 424350
rect 43274 424294 43342 424350
rect 43398 424294 43494 424350
rect 42874 424226 43494 424294
rect 42874 424170 42970 424226
rect 43026 424170 43094 424226
rect 43150 424170 43218 424226
rect 43274 424170 43342 424226
rect 43398 424170 43494 424226
rect 42874 424102 43494 424170
rect 42874 424046 42970 424102
rect 43026 424046 43094 424102
rect 43150 424046 43218 424102
rect 43274 424046 43342 424102
rect 43398 424046 43494 424102
rect 42874 423978 43494 424046
rect 42874 423922 42970 423978
rect 43026 423922 43094 423978
rect 43150 423922 43218 423978
rect 43274 423922 43342 423978
rect 43398 423922 43494 423978
rect 42874 406350 43494 423922
rect 54448 418350 54768 418384
rect 54448 418294 54518 418350
rect 54574 418294 54642 418350
rect 54698 418294 54768 418350
rect 54448 418226 54768 418294
rect 54448 418170 54518 418226
rect 54574 418170 54642 418226
rect 54698 418170 54768 418226
rect 54448 418102 54768 418170
rect 54448 418046 54518 418102
rect 54574 418046 54642 418102
rect 54698 418046 54768 418102
rect 54448 417978 54768 418046
rect 54448 417922 54518 417978
rect 54574 417922 54642 417978
rect 54698 417922 54768 417978
rect 54448 417888 54768 417922
rect 57154 418350 57774 435922
rect 57154 418294 57250 418350
rect 57306 418294 57374 418350
rect 57430 418294 57498 418350
rect 57554 418294 57622 418350
rect 57678 418294 57774 418350
rect 57154 418226 57774 418294
rect 57154 418170 57250 418226
rect 57306 418170 57374 418226
rect 57430 418170 57498 418226
rect 57554 418170 57622 418226
rect 57678 418170 57774 418226
rect 57154 418102 57774 418170
rect 57154 418046 57250 418102
rect 57306 418046 57374 418102
rect 57430 418046 57498 418102
rect 57554 418046 57622 418102
rect 57678 418046 57774 418102
rect 57154 417978 57774 418046
rect 57154 417922 57250 417978
rect 57306 417922 57374 417978
rect 57430 417922 57498 417978
rect 57554 417922 57622 417978
rect 57678 417922 57774 417978
rect 42874 406294 42970 406350
rect 43026 406294 43094 406350
rect 43150 406294 43218 406350
rect 43274 406294 43342 406350
rect 43398 406294 43494 406350
rect 42874 406226 43494 406294
rect 42874 406170 42970 406226
rect 43026 406170 43094 406226
rect 43150 406170 43218 406226
rect 43274 406170 43342 406226
rect 43398 406170 43494 406226
rect 42874 406102 43494 406170
rect 42874 406046 42970 406102
rect 43026 406046 43094 406102
rect 43150 406046 43218 406102
rect 43274 406046 43342 406102
rect 43398 406046 43494 406102
rect 42874 405978 43494 406046
rect 42874 405922 42970 405978
rect 43026 405922 43094 405978
rect 43150 405922 43218 405978
rect 43274 405922 43342 405978
rect 43398 405922 43494 405978
rect 42874 388350 43494 405922
rect 54448 400350 54768 400384
rect 54448 400294 54518 400350
rect 54574 400294 54642 400350
rect 54698 400294 54768 400350
rect 54448 400226 54768 400294
rect 54448 400170 54518 400226
rect 54574 400170 54642 400226
rect 54698 400170 54768 400226
rect 54448 400102 54768 400170
rect 54448 400046 54518 400102
rect 54574 400046 54642 400102
rect 54698 400046 54768 400102
rect 54448 399978 54768 400046
rect 54448 399922 54518 399978
rect 54574 399922 54642 399978
rect 54698 399922 54768 399978
rect 54448 399888 54768 399922
rect 57154 400350 57774 417922
rect 57154 400294 57250 400350
rect 57306 400294 57374 400350
rect 57430 400294 57498 400350
rect 57554 400294 57622 400350
rect 57678 400294 57774 400350
rect 57154 400226 57774 400294
rect 57154 400170 57250 400226
rect 57306 400170 57374 400226
rect 57430 400170 57498 400226
rect 57554 400170 57622 400226
rect 57678 400170 57774 400226
rect 57154 400102 57774 400170
rect 57154 400046 57250 400102
rect 57306 400046 57374 400102
rect 57430 400046 57498 400102
rect 57554 400046 57622 400102
rect 57678 400046 57774 400102
rect 57154 399978 57774 400046
rect 57154 399922 57250 399978
rect 57306 399922 57374 399978
rect 57430 399922 57498 399978
rect 57554 399922 57622 399978
rect 57678 399922 57774 399978
rect 42874 388294 42970 388350
rect 43026 388294 43094 388350
rect 43150 388294 43218 388350
rect 43274 388294 43342 388350
rect 43398 388294 43494 388350
rect 42874 388226 43494 388294
rect 42874 388170 42970 388226
rect 43026 388170 43094 388226
rect 43150 388170 43218 388226
rect 43274 388170 43342 388226
rect 43398 388170 43494 388226
rect 42874 388102 43494 388170
rect 42874 388046 42970 388102
rect 43026 388046 43094 388102
rect 43150 388046 43218 388102
rect 43274 388046 43342 388102
rect 43398 388046 43494 388102
rect 42874 387978 43494 388046
rect 42874 387922 42970 387978
rect 43026 387922 43094 387978
rect 43150 387922 43218 387978
rect 43274 387922 43342 387978
rect 43398 387922 43494 387978
rect 42874 370350 43494 387922
rect 54448 382350 54768 382384
rect 54448 382294 54518 382350
rect 54574 382294 54642 382350
rect 54698 382294 54768 382350
rect 54448 382226 54768 382294
rect 54448 382170 54518 382226
rect 54574 382170 54642 382226
rect 54698 382170 54768 382226
rect 54448 382102 54768 382170
rect 54448 382046 54518 382102
rect 54574 382046 54642 382102
rect 54698 382046 54768 382102
rect 54448 381978 54768 382046
rect 54448 381922 54518 381978
rect 54574 381922 54642 381978
rect 54698 381922 54768 381978
rect 54448 381888 54768 381922
rect 57154 382350 57774 399922
rect 57154 382294 57250 382350
rect 57306 382294 57374 382350
rect 57430 382294 57498 382350
rect 57554 382294 57622 382350
rect 57678 382294 57774 382350
rect 57154 382226 57774 382294
rect 57154 382170 57250 382226
rect 57306 382170 57374 382226
rect 57430 382170 57498 382226
rect 57554 382170 57622 382226
rect 57678 382170 57774 382226
rect 57154 382102 57774 382170
rect 57154 382046 57250 382102
rect 57306 382046 57374 382102
rect 57430 382046 57498 382102
rect 57554 382046 57622 382102
rect 57678 382046 57774 382102
rect 57154 381978 57774 382046
rect 57154 381922 57250 381978
rect 57306 381922 57374 381978
rect 57430 381922 57498 381978
rect 57554 381922 57622 381978
rect 57678 381922 57774 381978
rect 42874 370294 42970 370350
rect 43026 370294 43094 370350
rect 43150 370294 43218 370350
rect 43274 370294 43342 370350
rect 43398 370294 43494 370350
rect 42874 370226 43494 370294
rect 42874 370170 42970 370226
rect 43026 370170 43094 370226
rect 43150 370170 43218 370226
rect 43274 370170 43342 370226
rect 43398 370170 43494 370226
rect 42874 370102 43494 370170
rect 42874 370046 42970 370102
rect 43026 370046 43094 370102
rect 43150 370046 43218 370102
rect 43274 370046 43342 370102
rect 43398 370046 43494 370102
rect 42874 369978 43494 370046
rect 42874 369922 42970 369978
rect 43026 369922 43094 369978
rect 43150 369922 43218 369978
rect 43274 369922 43342 369978
rect 43398 369922 43494 369978
rect 42874 352350 43494 369922
rect 54448 364350 54768 364384
rect 54448 364294 54518 364350
rect 54574 364294 54642 364350
rect 54698 364294 54768 364350
rect 54448 364226 54768 364294
rect 54448 364170 54518 364226
rect 54574 364170 54642 364226
rect 54698 364170 54768 364226
rect 54448 364102 54768 364170
rect 54448 364046 54518 364102
rect 54574 364046 54642 364102
rect 54698 364046 54768 364102
rect 54448 363978 54768 364046
rect 54448 363922 54518 363978
rect 54574 363922 54642 363978
rect 54698 363922 54768 363978
rect 54448 363888 54768 363922
rect 57154 364350 57774 381922
rect 57154 364294 57250 364350
rect 57306 364294 57374 364350
rect 57430 364294 57498 364350
rect 57554 364294 57622 364350
rect 57678 364294 57774 364350
rect 57154 364226 57774 364294
rect 57154 364170 57250 364226
rect 57306 364170 57374 364226
rect 57430 364170 57498 364226
rect 57554 364170 57622 364226
rect 57678 364170 57774 364226
rect 57154 364102 57774 364170
rect 57154 364046 57250 364102
rect 57306 364046 57374 364102
rect 57430 364046 57498 364102
rect 57554 364046 57622 364102
rect 57678 364046 57774 364102
rect 57154 363978 57774 364046
rect 57154 363922 57250 363978
rect 57306 363922 57374 363978
rect 57430 363922 57498 363978
rect 57554 363922 57622 363978
rect 57678 363922 57774 363978
rect 42874 352294 42970 352350
rect 43026 352294 43094 352350
rect 43150 352294 43218 352350
rect 43274 352294 43342 352350
rect 43398 352294 43494 352350
rect 42874 352226 43494 352294
rect 42874 352170 42970 352226
rect 43026 352170 43094 352226
rect 43150 352170 43218 352226
rect 43274 352170 43342 352226
rect 43398 352170 43494 352226
rect 42874 352102 43494 352170
rect 42874 352046 42970 352102
rect 43026 352046 43094 352102
rect 43150 352046 43218 352102
rect 43274 352046 43342 352102
rect 43398 352046 43494 352102
rect 42874 351978 43494 352046
rect 42874 351922 42970 351978
rect 43026 351922 43094 351978
rect 43150 351922 43218 351978
rect 43274 351922 43342 351978
rect 43398 351922 43494 351978
rect 42874 334350 43494 351922
rect 54448 346350 54768 346384
rect 54448 346294 54518 346350
rect 54574 346294 54642 346350
rect 54698 346294 54768 346350
rect 54448 346226 54768 346294
rect 54448 346170 54518 346226
rect 54574 346170 54642 346226
rect 54698 346170 54768 346226
rect 54448 346102 54768 346170
rect 54448 346046 54518 346102
rect 54574 346046 54642 346102
rect 54698 346046 54768 346102
rect 54448 345978 54768 346046
rect 54448 345922 54518 345978
rect 54574 345922 54642 345978
rect 54698 345922 54768 345978
rect 54448 345888 54768 345922
rect 57154 346350 57774 363922
rect 57154 346294 57250 346350
rect 57306 346294 57374 346350
rect 57430 346294 57498 346350
rect 57554 346294 57622 346350
rect 57678 346294 57774 346350
rect 57154 346226 57774 346294
rect 57154 346170 57250 346226
rect 57306 346170 57374 346226
rect 57430 346170 57498 346226
rect 57554 346170 57622 346226
rect 57678 346170 57774 346226
rect 57154 346102 57774 346170
rect 57154 346046 57250 346102
rect 57306 346046 57374 346102
rect 57430 346046 57498 346102
rect 57554 346046 57622 346102
rect 57678 346046 57774 346102
rect 57154 345978 57774 346046
rect 57154 345922 57250 345978
rect 57306 345922 57374 345978
rect 57430 345922 57498 345978
rect 57554 345922 57622 345978
rect 57678 345922 57774 345978
rect 42874 334294 42970 334350
rect 43026 334294 43094 334350
rect 43150 334294 43218 334350
rect 43274 334294 43342 334350
rect 43398 334294 43494 334350
rect 42874 334226 43494 334294
rect 42874 334170 42970 334226
rect 43026 334170 43094 334226
rect 43150 334170 43218 334226
rect 43274 334170 43342 334226
rect 43398 334170 43494 334226
rect 42874 334102 43494 334170
rect 42874 334046 42970 334102
rect 43026 334046 43094 334102
rect 43150 334046 43218 334102
rect 43274 334046 43342 334102
rect 43398 334046 43494 334102
rect 42874 333978 43494 334046
rect 42874 333922 42970 333978
rect 43026 333922 43094 333978
rect 43150 333922 43218 333978
rect 43274 333922 43342 333978
rect 43398 333922 43494 333978
rect 42874 316350 43494 333922
rect 54448 328350 54768 328384
rect 54448 328294 54518 328350
rect 54574 328294 54642 328350
rect 54698 328294 54768 328350
rect 54448 328226 54768 328294
rect 54448 328170 54518 328226
rect 54574 328170 54642 328226
rect 54698 328170 54768 328226
rect 54448 328102 54768 328170
rect 54448 328046 54518 328102
rect 54574 328046 54642 328102
rect 54698 328046 54768 328102
rect 54448 327978 54768 328046
rect 54448 327922 54518 327978
rect 54574 327922 54642 327978
rect 54698 327922 54768 327978
rect 54448 327888 54768 327922
rect 57154 328350 57774 345922
rect 57154 328294 57250 328350
rect 57306 328294 57374 328350
rect 57430 328294 57498 328350
rect 57554 328294 57622 328350
rect 57678 328294 57774 328350
rect 57154 328226 57774 328294
rect 57154 328170 57250 328226
rect 57306 328170 57374 328226
rect 57430 328170 57498 328226
rect 57554 328170 57622 328226
rect 57678 328170 57774 328226
rect 57154 328102 57774 328170
rect 57154 328046 57250 328102
rect 57306 328046 57374 328102
rect 57430 328046 57498 328102
rect 57554 328046 57622 328102
rect 57678 328046 57774 328102
rect 57154 327978 57774 328046
rect 57154 327922 57250 327978
rect 57306 327922 57374 327978
rect 57430 327922 57498 327978
rect 57554 327922 57622 327978
rect 57678 327922 57774 327978
rect 42874 316294 42970 316350
rect 43026 316294 43094 316350
rect 43150 316294 43218 316350
rect 43274 316294 43342 316350
rect 43398 316294 43494 316350
rect 42874 316226 43494 316294
rect 42874 316170 42970 316226
rect 43026 316170 43094 316226
rect 43150 316170 43218 316226
rect 43274 316170 43342 316226
rect 43398 316170 43494 316226
rect 42874 316102 43494 316170
rect 42874 316046 42970 316102
rect 43026 316046 43094 316102
rect 43150 316046 43218 316102
rect 43274 316046 43342 316102
rect 43398 316046 43494 316102
rect 42874 315978 43494 316046
rect 42874 315922 42970 315978
rect 43026 315922 43094 315978
rect 43150 315922 43218 315978
rect 43274 315922 43342 315978
rect 43398 315922 43494 315978
rect 42874 298350 43494 315922
rect 54448 310350 54768 310384
rect 54448 310294 54518 310350
rect 54574 310294 54642 310350
rect 54698 310294 54768 310350
rect 54448 310226 54768 310294
rect 54448 310170 54518 310226
rect 54574 310170 54642 310226
rect 54698 310170 54768 310226
rect 54448 310102 54768 310170
rect 54448 310046 54518 310102
rect 54574 310046 54642 310102
rect 54698 310046 54768 310102
rect 54448 309978 54768 310046
rect 54448 309922 54518 309978
rect 54574 309922 54642 309978
rect 54698 309922 54768 309978
rect 54448 309888 54768 309922
rect 57154 310350 57774 327922
rect 57154 310294 57250 310350
rect 57306 310294 57374 310350
rect 57430 310294 57498 310350
rect 57554 310294 57622 310350
rect 57678 310294 57774 310350
rect 57154 310226 57774 310294
rect 57154 310170 57250 310226
rect 57306 310170 57374 310226
rect 57430 310170 57498 310226
rect 57554 310170 57622 310226
rect 57678 310170 57774 310226
rect 57154 310102 57774 310170
rect 57154 310046 57250 310102
rect 57306 310046 57374 310102
rect 57430 310046 57498 310102
rect 57554 310046 57622 310102
rect 57678 310046 57774 310102
rect 57154 309978 57774 310046
rect 57154 309922 57250 309978
rect 57306 309922 57374 309978
rect 57430 309922 57498 309978
rect 57554 309922 57622 309978
rect 57678 309922 57774 309978
rect 42874 298294 42970 298350
rect 43026 298294 43094 298350
rect 43150 298294 43218 298350
rect 43274 298294 43342 298350
rect 43398 298294 43494 298350
rect 42874 298226 43494 298294
rect 42874 298170 42970 298226
rect 43026 298170 43094 298226
rect 43150 298170 43218 298226
rect 43274 298170 43342 298226
rect 43398 298170 43494 298226
rect 42874 298102 43494 298170
rect 42874 298046 42970 298102
rect 43026 298046 43094 298102
rect 43150 298046 43218 298102
rect 43274 298046 43342 298102
rect 43398 298046 43494 298102
rect 42874 297978 43494 298046
rect 42874 297922 42970 297978
rect 43026 297922 43094 297978
rect 43150 297922 43218 297978
rect 43274 297922 43342 297978
rect 43398 297922 43494 297978
rect 42874 280350 43494 297922
rect 54448 292350 54768 292384
rect 54448 292294 54518 292350
rect 54574 292294 54642 292350
rect 54698 292294 54768 292350
rect 54448 292226 54768 292294
rect 54448 292170 54518 292226
rect 54574 292170 54642 292226
rect 54698 292170 54768 292226
rect 54448 292102 54768 292170
rect 54448 292046 54518 292102
rect 54574 292046 54642 292102
rect 54698 292046 54768 292102
rect 54448 291978 54768 292046
rect 54448 291922 54518 291978
rect 54574 291922 54642 291978
rect 54698 291922 54768 291978
rect 54448 291888 54768 291922
rect 57154 292350 57774 309922
rect 57154 292294 57250 292350
rect 57306 292294 57374 292350
rect 57430 292294 57498 292350
rect 57554 292294 57622 292350
rect 57678 292294 57774 292350
rect 57154 292226 57774 292294
rect 57154 292170 57250 292226
rect 57306 292170 57374 292226
rect 57430 292170 57498 292226
rect 57554 292170 57622 292226
rect 57678 292170 57774 292226
rect 57154 292102 57774 292170
rect 57154 292046 57250 292102
rect 57306 292046 57374 292102
rect 57430 292046 57498 292102
rect 57554 292046 57622 292102
rect 57678 292046 57774 292102
rect 57154 291978 57774 292046
rect 57154 291922 57250 291978
rect 57306 291922 57374 291978
rect 57430 291922 57498 291978
rect 57554 291922 57622 291978
rect 57678 291922 57774 291978
rect 42874 280294 42970 280350
rect 43026 280294 43094 280350
rect 43150 280294 43218 280350
rect 43274 280294 43342 280350
rect 43398 280294 43494 280350
rect 42874 280226 43494 280294
rect 42874 280170 42970 280226
rect 43026 280170 43094 280226
rect 43150 280170 43218 280226
rect 43274 280170 43342 280226
rect 43398 280170 43494 280226
rect 42874 280102 43494 280170
rect 42874 280046 42970 280102
rect 43026 280046 43094 280102
rect 43150 280046 43218 280102
rect 43274 280046 43342 280102
rect 43398 280046 43494 280102
rect 42874 279978 43494 280046
rect 42874 279922 42970 279978
rect 43026 279922 43094 279978
rect 43150 279922 43218 279978
rect 43274 279922 43342 279978
rect 43398 279922 43494 279978
rect 42874 262350 43494 279922
rect 54448 274350 54768 274384
rect 54448 274294 54518 274350
rect 54574 274294 54642 274350
rect 54698 274294 54768 274350
rect 54448 274226 54768 274294
rect 54448 274170 54518 274226
rect 54574 274170 54642 274226
rect 54698 274170 54768 274226
rect 54448 274102 54768 274170
rect 54448 274046 54518 274102
rect 54574 274046 54642 274102
rect 54698 274046 54768 274102
rect 54448 273978 54768 274046
rect 54448 273922 54518 273978
rect 54574 273922 54642 273978
rect 54698 273922 54768 273978
rect 54448 273888 54768 273922
rect 57154 274350 57774 291922
rect 57154 274294 57250 274350
rect 57306 274294 57374 274350
rect 57430 274294 57498 274350
rect 57554 274294 57622 274350
rect 57678 274294 57774 274350
rect 57154 274226 57774 274294
rect 57154 274170 57250 274226
rect 57306 274170 57374 274226
rect 57430 274170 57498 274226
rect 57554 274170 57622 274226
rect 57678 274170 57774 274226
rect 57154 274102 57774 274170
rect 57154 274046 57250 274102
rect 57306 274046 57374 274102
rect 57430 274046 57498 274102
rect 57554 274046 57622 274102
rect 57678 274046 57774 274102
rect 57154 273978 57774 274046
rect 57154 273922 57250 273978
rect 57306 273922 57374 273978
rect 57430 273922 57498 273978
rect 57554 273922 57622 273978
rect 57678 273922 57774 273978
rect 42874 262294 42970 262350
rect 43026 262294 43094 262350
rect 43150 262294 43218 262350
rect 43274 262294 43342 262350
rect 43398 262294 43494 262350
rect 42874 262226 43494 262294
rect 42874 262170 42970 262226
rect 43026 262170 43094 262226
rect 43150 262170 43218 262226
rect 43274 262170 43342 262226
rect 43398 262170 43494 262226
rect 42874 262102 43494 262170
rect 42874 262046 42970 262102
rect 43026 262046 43094 262102
rect 43150 262046 43218 262102
rect 43274 262046 43342 262102
rect 43398 262046 43494 262102
rect 42874 261978 43494 262046
rect 42874 261922 42970 261978
rect 43026 261922 43094 261978
rect 43150 261922 43218 261978
rect 43274 261922 43342 261978
rect 43398 261922 43494 261978
rect 42874 244350 43494 261922
rect 54448 256350 54768 256384
rect 54448 256294 54518 256350
rect 54574 256294 54642 256350
rect 54698 256294 54768 256350
rect 54448 256226 54768 256294
rect 54448 256170 54518 256226
rect 54574 256170 54642 256226
rect 54698 256170 54768 256226
rect 54448 256102 54768 256170
rect 54448 256046 54518 256102
rect 54574 256046 54642 256102
rect 54698 256046 54768 256102
rect 54448 255978 54768 256046
rect 54448 255922 54518 255978
rect 54574 255922 54642 255978
rect 54698 255922 54768 255978
rect 54448 255888 54768 255922
rect 57154 256350 57774 273922
rect 57154 256294 57250 256350
rect 57306 256294 57374 256350
rect 57430 256294 57498 256350
rect 57554 256294 57622 256350
rect 57678 256294 57774 256350
rect 57154 256226 57774 256294
rect 57154 256170 57250 256226
rect 57306 256170 57374 256226
rect 57430 256170 57498 256226
rect 57554 256170 57622 256226
rect 57678 256170 57774 256226
rect 57154 256102 57774 256170
rect 57154 256046 57250 256102
rect 57306 256046 57374 256102
rect 57430 256046 57498 256102
rect 57554 256046 57622 256102
rect 57678 256046 57774 256102
rect 57154 255978 57774 256046
rect 57154 255922 57250 255978
rect 57306 255922 57374 255978
rect 57430 255922 57498 255978
rect 57554 255922 57622 255978
rect 57678 255922 57774 255978
rect 42874 244294 42970 244350
rect 43026 244294 43094 244350
rect 43150 244294 43218 244350
rect 43274 244294 43342 244350
rect 43398 244294 43494 244350
rect 42874 244226 43494 244294
rect 42874 244170 42970 244226
rect 43026 244170 43094 244226
rect 43150 244170 43218 244226
rect 43274 244170 43342 244226
rect 43398 244170 43494 244226
rect 42874 244102 43494 244170
rect 42874 244046 42970 244102
rect 43026 244046 43094 244102
rect 43150 244046 43218 244102
rect 43274 244046 43342 244102
rect 43398 244046 43494 244102
rect 42874 243978 43494 244046
rect 42874 243922 42970 243978
rect 43026 243922 43094 243978
rect 43150 243922 43218 243978
rect 43274 243922 43342 243978
rect 43398 243922 43494 243978
rect 42874 226350 43494 243922
rect 54448 238350 54768 238384
rect 54448 238294 54518 238350
rect 54574 238294 54642 238350
rect 54698 238294 54768 238350
rect 54448 238226 54768 238294
rect 54448 238170 54518 238226
rect 54574 238170 54642 238226
rect 54698 238170 54768 238226
rect 54448 238102 54768 238170
rect 54448 238046 54518 238102
rect 54574 238046 54642 238102
rect 54698 238046 54768 238102
rect 54448 237978 54768 238046
rect 54448 237922 54518 237978
rect 54574 237922 54642 237978
rect 54698 237922 54768 237978
rect 54448 237888 54768 237922
rect 57154 238350 57774 255922
rect 57154 238294 57250 238350
rect 57306 238294 57374 238350
rect 57430 238294 57498 238350
rect 57554 238294 57622 238350
rect 57678 238294 57774 238350
rect 57154 238226 57774 238294
rect 57154 238170 57250 238226
rect 57306 238170 57374 238226
rect 57430 238170 57498 238226
rect 57554 238170 57622 238226
rect 57678 238170 57774 238226
rect 57154 238102 57774 238170
rect 57154 238046 57250 238102
rect 57306 238046 57374 238102
rect 57430 238046 57498 238102
rect 57554 238046 57622 238102
rect 57678 238046 57774 238102
rect 57154 237978 57774 238046
rect 57154 237922 57250 237978
rect 57306 237922 57374 237978
rect 57430 237922 57498 237978
rect 57554 237922 57622 237978
rect 57678 237922 57774 237978
rect 49868 237748 49924 237758
rect 50204 237748 50260 237758
rect 49924 237692 50204 237748
rect 49868 237682 49924 237692
rect 50204 237682 50260 237692
rect 42874 226294 42970 226350
rect 43026 226294 43094 226350
rect 43150 226294 43218 226350
rect 43274 226294 43342 226350
rect 43398 226294 43494 226350
rect 42874 226226 43494 226294
rect 42874 226170 42970 226226
rect 43026 226170 43094 226226
rect 43150 226170 43218 226226
rect 43274 226170 43342 226226
rect 43398 226170 43494 226226
rect 42874 226102 43494 226170
rect 42874 226046 42970 226102
rect 43026 226046 43094 226102
rect 43150 226046 43218 226102
rect 43274 226046 43342 226102
rect 43398 226046 43494 226102
rect 42874 225978 43494 226046
rect 42874 225922 42970 225978
rect 43026 225922 43094 225978
rect 43150 225922 43218 225978
rect 43274 225922 43342 225978
rect 43398 225922 43494 225978
rect 42874 208350 43494 225922
rect 54448 220350 54768 220384
rect 54448 220294 54518 220350
rect 54574 220294 54642 220350
rect 54698 220294 54768 220350
rect 54448 220226 54768 220294
rect 54448 220170 54518 220226
rect 54574 220170 54642 220226
rect 54698 220170 54768 220226
rect 54448 220102 54768 220170
rect 54448 220046 54518 220102
rect 54574 220046 54642 220102
rect 54698 220046 54768 220102
rect 54448 219978 54768 220046
rect 54448 219922 54518 219978
rect 54574 219922 54642 219978
rect 54698 219922 54768 219978
rect 54448 219888 54768 219922
rect 57154 220350 57774 237922
rect 57154 220294 57250 220350
rect 57306 220294 57374 220350
rect 57430 220294 57498 220350
rect 57554 220294 57622 220350
rect 57678 220294 57774 220350
rect 57154 220226 57774 220294
rect 57154 220170 57250 220226
rect 57306 220170 57374 220226
rect 57430 220170 57498 220226
rect 57554 220170 57622 220226
rect 57678 220170 57774 220226
rect 57154 220102 57774 220170
rect 57154 220046 57250 220102
rect 57306 220046 57374 220102
rect 57430 220046 57498 220102
rect 57554 220046 57622 220102
rect 57678 220046 57774 220102
rect 57154 219978 57774 220046
rect 57154 219922 57250 219978
rect 57306 219922 57374 219978
rect 57430 219922 57498 219978
rect 57554 219922 57622 219978
rect 57678 219922 57774 219978
rect 42874 208294 42970 208350
rect 43026 208294 43094 208350
rect 43150 208294 43218 208350
rect 43274 208294 43342 208350
rect 43398 208294 43494 208350
rect 42874 208226 43494 208294
rect 42874 208170 42970 208226
rect 43026 208170 43094 208226
rect 43150 208170 43218 208226
rect 43274 208170 43342 208226
rect 43398 208170 43494 208226
rect 42874 208102 43494 208170
rect 42874 208046 42970 208102
rect 43026 208046 43094 208102
rect 43150 208046 43218 208102
rect 43274 208046 43342 208102
rect 43398 208046 43494 208102
rect 42874 207978 43494 208046
rect 42874 207922 42970 207978
rect 43026 207922 43094 207978
rect 43150 207922 43218 207978
rect 43274 207922 43342 207978
rect 43398 207922 43494 207978
rect 42874 190350 43494 207922
rect 54448 202350 54768 202384
rect 54448 202294 54518 202350
rect 54574 202294 54642 202350
rect 54698 202294 54768 202350
rect 54448 202226 54768 202294
rect 54448 202170 54518 202226
rect 54574 202170 54642 202226
rect 54698 202170 54768 202226
rect 54448 202102 54768 202170
rect 54448 202046 54518 202102
rect 54574 202046 54642 202102
rect 54698 202046 54768 202102
rect 54448 201978 54768 202046
rect 54448 201922 54518 201978
rect 54574 201922 54642 201978
rect 54698 201922 54768 201978
rect 54448 201888 54768 201922
rect 57154 202350 57774 219922
rect 57154 202294 57250 202350
rect 57306 202294 57374 202350
rect 57430 202294 57498 202350
rect 57554 202294 57622 202350
rect 57678 202294 57774 202350
rect 57154 202226 57774 202294
rect 57154 202170 57250 202226
rect 57306 202170 57374 202226
rect 57430 202170 57498 202226
rect 57554 202170 57622 202226
rect 57678 202170 57774 202226
rect 57154 202102 57774 202170
rect 57154 202046 57250 202102
rect 57306 202046 57374 202102
rect 57430 202046 57498 202102
rect 57554 202046 57622 202102
rect 57678 202046 57774 202102
rect 57154 201978 57774 202046
rect 57154 201922 57250 201978
rect 57306 201922 57374 201978
rect 57430 201922 57498 201978
rect 57554 201922 57622 201978
rect 57678 201922 57774 201978
rect 42874 190294 42970 190350
rect 43026 190294 43094 190350
rect 43150 190294 43218 190350
rect 43274 190294 43342 190350
rect 43398 190294 43494 190350
rect 42874 190226 43494 190294
rect 42874 190170 42970 190226
rect 43026 190170 43094 190226
rect 43150 190170 43218 190226
rect 43274 190170 43342 190226
rect 43398 190170 43494 190226
rect 42874 190102 43494 190170
rect 42874 190046 42970 190102
rect 43026 190046 43094 190102
rect 43150 190046 43218 190102
rect 43274 190046 43342 190102
rect 43398 190046 43494 190102
rect 42874 189978 43494 190046
rect 42874 189922 42970 189978
rect 43026 189922 43094 189978
rect 43150 189922 43218 189978
rect 43274 189922 43342 189978
rect 43398 189922 43494 189978
rect 42874 172350 43494 189922
rect 54448 184350 54768 184384
rect 54448 184294 54518 184350
rect 54574 184294 54642 184350
rect 54698 184294 54768 184350
rect 54448 184226 54768 184294
rect 54448 184170 54518 184226
rect 54574 184170 54642 184226
rect 54698 184170 54768 184226
rect 54448 184102 54768 184170
rect 54448 184046 54518 184102
rect 54574 184046 54642 184102
rect 54698 184046 54768 184102
rect 54448 183978 54768 184046
rect 54448 183922 54518 183978
rect 54574 183922 54642 183978
rect 54698 183922 54768 183978
rect 54448 183888 54768 183922
rect 57154 184350 57774 201922
rect 57154 184294 57250 184350
rect 57306 184294 57374 184350
rect 57430 184294 57498 184350
rect 57554 184294 57622 184350
rect 57678 184294 57774 184350
rect 57154 184226 57774 184294
rect 57154 184170 57250 184226
rect 57306 184170 57374 184226
rect 57430 184170 57498 184226
rect 57554 184170 57622 184226
rect 57678 184170 57774 184226
rect 57154 184102 57774 184170
rect 57154 184046 57250 184102
rect 57306 184046 57374 184102
rect 57430 184046 57498 184102
rect 57554 184046 57622 184102
rect 57678 184046 57774 184102
rect 57154 183978 57774 184046
rect 57154 183922 57250 183978
rect 57306 183922 57374 183978
rect 57430 183922 57498 183978
rect 57554 183922 57622 183978
rect 57678 183922 57774 183978
rect 42874 172294 42970 172350
rect 43026 172294 43094 172350
rect 43150 172294 43218 172350
rect 43274 172294 43342 172350
rect 43398 172294 43494 172350
rect 42874 172226 43494 172294
rect 42874 172170 42970 172226
rect 43026 172170 43094 172226
rect 43150 172170 43218 172226
rect 43274 172170 43342 172226
rect 43398 172170 43494 172226
rect 42874 172102 43494 172170
rect 42874 172046 42970 172102
rect 43026 172046 43094 172102
rect 43150 172046 43218 172102
rect 43274 172046 43342 172102
rect 43398 172046 43494 172102
rect 42874 171978 43494 172046
rect 42874 171922 42970 171978
rect 43026 171922 43094 171978
rect 43150 171922 43218 171978
rect 43274 171922 43342 171978
rect 43398 171922 43494 171978
rect 42874 154350 43494 171922
rect 54448 166350 54768 166384
rect 54448 166294 54518 166350
rect 54574 166294 54642 166350
rect 54698 166294 54768 166350
rect 54448 166226 54768 166294
rect 54448 166170 54518 166226
rect 54574 166170 54642 166226
rect 54698 166170 54768 166226
rect 54448 166102 54768 166170
rect 54448 166046 54518 166102
rect 54574 166046 54642 166102
rect 54698 166046 54768 166102
rect 54448 165978 54768 166046
rect 54448 165922 54518 165978
rect 54574 165922 54642 165978
rect 54698 165922 54768 165978
rect 54448 165888 54768 165922
rect 57154 166350 57774 183922
rect 57154 166294 57250 166350
rect 57306 166294 57374 166350
rect 57430 166294 57498 166350
rect 57554 166294 57622 166350
rect 57678 166294 57774 166350
rect 57154 166226 57774 166294
rect 57154 166170 57250 166226
rect 57306 166170 57374 166226
rect 57430 166170 57498 166226
rect 57554 166170 57622 166226
rect 57678 166170 57774 166226
rect 57154 166102 57774 166170
rect 57154 166046 57250 166102
rect 57306 166046 57374 166102
rect 57430 166046 57498 166102
rect 57554 166046 57622 166102
rect 57678 166046 57774 166102
rect 57154 165978 57774 166046
rect 57154 165922 57250 165978
rect 57306 165922 57374 165978
rect 57430 165922 57498 165978
rect 57554 165922 57622 165978
rect 57678 165922 57774 165978
rect 42874 154294 42970 154350
rect 43026 154294 43094 154350
rect 43150 154294 43218 154350
rect 43274 154294 43342 154350
rect 43398 154294 43494 154350
rect 42874 154226 43494 154294
rect 42874 154170 42970 154226
rect 43026 154170 43094 154226
rect 43150 154170 43218 154226
rect 43274 154170 43342 154226
rect 43398 154170 43494 154226
rect 42874 154102 43494 154170
rect 42874 154046 42970 154102
rect 43026 154046 43094 154102
rect 43150 154046 43218 154102
rect 43274 154046 43342 154102
rect 43398 154046 43494 154102
rect 42874 153978 43494 154046
rect 42874 153922 42970 153978
rect 43026 153922 43094 153978
rect 43150 153922 43218 153978
rect 43274 153922 43342 153978
rect 43398 153922 43494 153978
rect 42874 136350 43494 153922
rect 54448 148350 54768 148384
rect 54448 148294 54518 148350
rect 54574 148294 54642 148350
rect 54698 148294 54768 148350
rect 54448 148226 54768 148294
rect 54448 148170 54518 148226
rect 54574 148170 54642 148226
rect 54698 148170 54768 148226
rect 54448 148102 54768 148170
rect 54448 148046 54518 148102
rect 54574 148046 54642 148102
rect 54698 148046 54768 148102
rect 54448 147978 54768 148046
rect 54448 147922 54518 147978
rect 54574 147922 54642 147978
rect 54698 147922 54768 147978
rect 54448 147888 54768 147922
rect 57154 148350 57774 165922
rect 57154 148294 57250 148350
rect 57306 148294 57374 148350
rect 57430 148294 57498 148350
rect 57554 148294 57622 148350
rect 57678 148294 57774 148350
rect 57154 148226 57774 148294
rect 57154 148170 57250 148226
rect 57306 148170 57374 148226
rect 57430 148170 57498 148226
rect 57554 148170 57622 148226
rect 57678 148170 57774 148226
rect 57154 148102 57774 148170
rect 57154 148046 57250 148102
rect 57306 148046 57374 148102
rect 57430 148046 57498 148102
rect 57554 148046 57622 148102
rect 57678 148046 57774 148102
rect 57154 147978 57774 148046
rect 57154 147922 57250 147978
rect 57306 147922 57374 147978
rect 57430 147922 57498 147978
rect 57554 147922 57622 147978
rect 57678 147922 57774 147978
rect 42874 136294 42970 136350
rect 43026 136294 43094 136350
rect 43150 136294 43218 136350
rect 43274 136294 43342 136350
rect 43398 136294 43494 136350
rect 42874 136226 43494 136294
rect 42874 136170 42970 136226
rect 43026 136170 43094 136226
rect 43150 136170 43218 136226
rect 43274 136170 43342 136226
rect 43398 136170 43494 136226
rect 42874 136102 43494 136170
rect 42874 136046 42970 136102
rect 43026 136046 43094 136102
rect 43150 136046 43218 136102
rect 43274 136046 43342 136102
rect 43398 136046 43494 136102
rect 42874 135978 43494 136046
rect 42874 135922 42970 135978
rect 43026 135922 43094 135978
rect 43150 135922 43218 135978
rect 43274 135922 43342 135978
rect 43398 135922 43494 135978
rect 42874 118350 43494 135922
rect 54448 130350 54768 130384
rect 54448 130294 54518 130350
rect 54574 130294 54642 130350
rect 54698 130294 54768 130350
rect 54448 130226 54768 130294
rect 54448 130170 54518 130226
rect 54574 130170 54642 130226
rect 54698 130170 54768 130226
rect 54448 130102 54768 130170
rect 54448 130046 54518 130102
rect 54574 130046 54642 130102
rect 54698 130046 54768 130102
rect 54448 129978 54768 130046
rect 54448 129922 54518 129978
rect 54574 129922 54642 129978
rect 54698 129922 54768 129978
rect 54448 129888 54768 129922
rect 57154 130350 57774 147922
rect 57154 130294 57250 130350
rect 57306 130294 57374 130350
rect 57430 130294 57498 130350
rect 57554 130294 57622 130350
rect 57678 130294 57774 130350
rect 57154 130226 57774 130294
rect 57154 130170 57250 130226
rect 57306 130170 57374 130226
rect 57430 130170 57498 130226
rect 57554 130170 57622 130226
rect 57678 130170 57774 130226
rect 57154 130102 57774 130170
rect 57154 130046 57250 130102
rect 57306 130046 57374 130102
rect 57430 130046 57498 130102
rect 57554 130046 57622 130102
rect 57678 130046 57774 130102
rect 57154 129978 57774 130046
rect 57154 129922 57250 129978
rect 57306 129922 57374 129978
rect 57430 129922 57498 129978
rect 57554 129922 57622 129978
rect 57678 129922 57774 129978
rect 42874 118294 42970 118350
rect 43026 118294 43094 118350
rect 43150 118294 43218 118350
rect 43274 118294 43342 118350
rect 43398 118294 43494 118350
rect 42874 118226 43494 118294
rect 42874 118170 42970 118226
rect 43026 118170 43094 118226
rect 43150 118170 43218 118226
rect 43274 118170 43342 118226
rect 43398 118170 43494 118226
rect 42874 118102 43494 118170
rect 42874 118046 42970 118102
rect 43026 118046 43094 118102
rect 43150 118046 43218 118102
rect 43274 118046 43342 118102
rect 43398 118046 43494 118102
rect 42874 117978 43494 118046
rect 42874 117922 42970 117978
rect 43026 117922 43094 117978
rect 43150 117922 43218 117978
rect 43274 117922 43342 117978
rect 43398 117922 43494 117978
rect 42874 100350 43494 117922
rect 54448 112350 54768 112384
rect 54448 112294 54518 112350
rect 54574 112294 54642 112350
rect 54698 112294 54768 112350
rect 54448 112226 54768 112294
rect 54448 112170 54518 112226
rect 54574 112170 54642 112226
rect 54698 112170 54768 112226
rect 54448 112102 54768 112170
rect 54448 112046 54518 112102
rect 54574 112046 54642 112102
rect 54698 112046 54768 112102
rect 54448 111978 54768 112046
rect 54448 111922 54518 111978
rect 54574 111922 54642 111978
rect 54698 111922 54768 111978
rect 54448 111888 54768 111922
rect 57154 112350 57774 129922
rect 57154 112294 57250 112350
rect 57306 112294 57374 112350
rect 57430 112294 57498 112350
rect 57554 112294 57622 112350
rect 57678 112294 57774 112350
rect 57154 112226 57774 112294
rect 57154 112170 57250 112226
rect 57306 112170 57374 112226
rect 57430 112170 57498 112226
rect 57554 112170 57622 112226
rect 57678 112170 57774 112226
rect 57154 112102 57774 112170
rect 57154 112046 57250 112102
rect 57306 112046 57374 112102
rect 57430 112046 57498 112102
rect 57554 112046 57622 112102
rect 57678 112046 57774 112102
rect 57154 111978 57774 112046
rect 57154 111922 57250 111978
rect 57306 111922 57374 111978
rect 57430 111922 57498 111978
rect 57554 111922 57622 111978
rect 57678 111922 57774 111978
rect 42874 100294 42970 100350
rect 43026 100294 43094 100350
rect 43150 100294 43218 100350
rect 43274 100294 43342 100350
rect 43398 100294 43494 100350
rect 42874 100226 43494 100294
rect 42874 100170 42970 100226
rect 43026 100170 43094 100226
rect 43150 100170 43218 100226
rect 43274 100170 43342 100226
rect 43398 100170 43494 100226
rect 42874 100102 43494 100170
rect 42874 100046 42970 100102
rect 43026 100046 43094 100102
rect 43150 100046 43218 100102
rect 43274 100046 43342 100102
rect 43398 100046 43494 100102
rect 42874 99978 43494 100046
rect 42874 99922 42970 99978
rect 43026 99922 43094 99978
rect 43150 99922 43218 99978
rect 43274 99922 43342 99978
rect 43398 99922 43494 99978
rect 42874 82350 43494 99922
rect 54448 94350 54768 94384
rect 54448 94294 54518 94350
rect 54574 94294 54642 94350
rect 54698 94294 54768 94350
rect 54448 94226 54768 94294
rect 54448 94170 54518 94226
rect 54574 94170 54642 94226
rect 54698 94170 54768 94226
rect 54448 94102 54768 94170
rect 54448 94046 54518 94102
rect 54574 94046 54642 94102
rect 54698 94046 54768 94102
rect 54448 93978 54768 94046
rect 54448 93922 54518 93978
rect 54574 93922 54642 93978
rect 54698 93922 54768 93978
rect 54448 93888 54768 93922
rect 57154 94350 57774 111922
rect 57154 94294 57250 94350
rect 57306 94294 57374 94350
rect 57430 94294 57498 94350
rect 57554 94294 57622 94350
rect 57678 94294 57774 94350
rect 57154 94226 57774 94294
rect 57154 94170 57250 94226
rect 57306 94170 57374 94226
rect 57430 94170 57498 94226
rect 57554 94170 57622 94226
rect 57678 94170 57774 94226
rect 57154 94102 57774 94170
rect 57154 94046 57250 94102
rect 57306 94046 57374 94102
rect 57430 94046 57498 94102
rect 57554 94046 57622 94102
rect 57678 94046 57774 94102
rect 57154 93978 57774 94046
rect 57154 93922 57250 93978
rect 57306 93922 57374 93978
rect 57430 93922 57498 93978
rect 57554 93922 57622 93978
rect 57678 93922 57774 93978
rect 42874 82294 42970 82350
rect 43026 82294 43094 82350
rect 43150 82294 43218 82350
rect 43274 82294 43342 82350
rect 43398 82294 43494 82350
rect 42874 82226 43494 82294
rect 42874 82170 42970 82226
rect 43026 82170 43094 82226
rect 43150 82170 43218 82226
rect 43274 82170 43342 82226
rect 43398 82170 43494 82226
rect 42874 82102 43494 82170
rect 42874 82046 42970 82102
rect 43026 82046 43094 82102
rect 43150 82046 43218 82102
rect 43274 82046 43342 82102
rect 43398 82046 43494 82102
rect 42874 81978 43494 82046
rect 42874 81922 42970 81978
rect 43026 81922 43094 81978
rect 43150 81922 43218 81978
rect 43274 81922 43342 81978
rect 43398 81922 43494 81978
rect 42874 64350 43494 81922
rect 54448 76350 54768 76384
rect 54448 76294 54518 76350
rect 54574 76294 54642 76350
rect 54698 76294 54768 76350
rect 54448 76226 54768 76294
rect 54448 76170 54518 76226
rect 54574 76170 54642 76226
rect 54698 76170 54768 76226
rect 54448 76102 54768 76170
rect 54448 76046 54518 76102
rect 54574 76046 54642 76102
rect 54698 76046 54768 76102
rect 54448 75978 54768 76046
rect 54448 75922 54518 75978
rect 54574 75922 54642 75978
rect 54698 75922 54768 75978
rect 54448 75888 54768 75922
rect 57154 76350 57774 93922
rect 57154 76294 57250 76350
rect 57306 76294 57374 76350
rect 57430 76294 57498 76350
rect 57554 76294 57622 76350
rect 57678 76294 57774 76350
rect 57154 76226 57774 76294
rect 57154 76170 57250 76226
rect 57306 76170 57374 76226
rect 57430 76170 57498 76226
rect 57554 76170 57622 76226
rect 57678 76170 57774 76226
rect 57154 76102 57774 76170
rect 57154 76046 57250 76102
rect 57306 76046 57374 76102
rect 57430 76046 57498 76102
rect 57554 76046 57622 76102
rect 57678 76046 57774 76102
rect 57154 75978 57774 76046
rect 57154 75922 57250 75978
rect 57306 75922 57374 75978
rect 57430 75922 57498 75978
rect 57554 75922 57622 75978
rect 57678 75922 57774 75978
rect 42874 64294 42970 64350
rect 43026 64294 43094 64350
rect 43150 64294 43218 64350
rect 43274 64294 43342 64350
rect 43398 64294 43494 64350
rect 42874 64226 43494 64294
rect 42874 64170 42970 64226
rect 43026 64170 43094 64226
rect 43150 64170 43218 64226
rect 43274 64170 43342 64226
rect 43398 64170 43494 64226
rect 42874 64102 43494 64170
rect 42874 64046 42970 64102
rect 43026 64046 43094 64102
rect 43150 64046 43218 64102
rect 43274 64046 43342 64102
rect 43398 64046 43494 64102
rect 42874 63978 43494 64046
rect 42874 63922 42970 63978
rect 43026 63922 43094 63978
rect 43150 63922 43218 63978
rect 43274 63922 43342 63978
rect 43398 63922 43494 63978
rect 42874 46350 43494 63922
rect 54448 58350 54768 58384
rect 54448 58294 54518 58350
rect 54574 58294 54642 58350
rect 54698 58294 54768 58350
rect 54448 58226 54768 58294
rect 54448 58170 54518 58226
rect 54574 58170 54642 58226
rect 54698 58170 54768 58226
rect 54448 58102 54768 58170
rect 54448 58046 54518 58102
rect 54574 58046 54642 58102
rect 54698 58046 54768 58102
rect 54448 57978 54768 58046
rect 54448 57922 54518 57978
rect 54574 57922 54642 57978
rect 54698 57922 54768 57978
rect 54448 57888 54768 57922
rect 57154 58350 57774 75922
rect 57154 58294 57250 58350
rect 57306 58294 57374 58350
rect 57430 58294 57498 58350
rect 57554 58294 57622 58350
rect 57678 58294 57774 58350
rect 57154 58226 57774 58294
rect 57154 58170 57250 58226
rect 57306 58170 57374 58226
rect 57430 58170 57498 58226
rect 57554 58170 57622 58226
rect 57678 58170 57774 58226
rect 57154 58102 57774 58170
rect 57154 58046 57250 58102
rect 57306 58046 57374 58102
rect 57430 58046 57498 58102
rect 57554 58046 57622 58102
rect 57678 58046 57774 58102
rect 57154 57978 57774 58046
rect 57154 57922 57250 57978
rect 57306 57922 57374 57978
rect 57430 57922 57498 57978
rect 57554 57922 57622 57978
rect 57678 57922 57774 57978
rect 42874 46294 42970 46350
rect 43026 46294 43094 46350
rect 43150 46294 43218 46350
rect 43274 46294 43342 46350
rect 43398 46294 43494 46350
rect 42874 46226 43494 46294
rect 42874 46170 42970 46226
rect 43026 46170 43094 46226
rect 43150 46170 43218 46226
rect 43274 46170 43342 46226
rect 43398 46170 43494 46226
rect 42874 46102 43494 46170
rect 42874 46046 42970 46102
rect 43026 46046 43094 46102
rect 43150 46046 43218 46102
rect 43274 46046 43342 46102
rect 43398 46046 43494 46102
rect 42874 45978 43494 46046
rect 42874 45922 42970 45978
rect 43026 45922 43094 45978
rect 43150 45922 43218 45978
rect 43274 45922 43342 45978
rect 43398 45922 43494 45978
rect 42874 28350 43494 45922
rect 54448 40350 54768 40384
rect 54448 40294 54518 40350
rect 54574 40294 54642 40350
rect 54698 40294 54768 40350
rect 54448 40226 54768 40294
rect 54448 40170 54518 40226
rect 54574 40170 54642 40226
rect 54698 40170 54768 40226
rect 54448 40102 54768 40170
rect 54448 40046 54518 40102
rect 54574 40046 54642 40102
rect 54698 40046 54768 40102
rect 54448 39978 54768 40046
rect 54448 39922 54518 39978
rect 54574 39922 54642 39978
rect 54698 39922 54768 39978
rect 54448 39888 54768 39922
rect 57154 40350 57774 57922
rect 57154 40294 57250 40350
rect 57306 40294 57374 40350
rect 57430 40294 57498 40350
rect 57554 40294 57622 40350
rect 57678 40294 57774 40350
rect 57154 40226 57774 40294
rect 57154 40170 57250 40226
rect 57306 40170 57374 40226
rect 57430 40170 57498 40226
rect 57554 40170 57622 40226
rect 57678 40170 57774 40226
rect 57154 40102 57774 40170
rect 57154 40046 57250 40102
rect 57306 40046 57374 40102
rect 57430 40046 57498 40102
rect 57554 40046 57622 40102
rect 57678 40046 57774 40102
rect 57154 39978 57774 40046
rect 57154 39922 57250 39978
rect 57306 39922 57374 39978
rect 57430 39922 57498 39978
rect 57554 39922 57622 39978
rect 57678 39922 57774 39978
rect 42874 28294 42970 28350
rect 43026 28294 43094 28350
rect 43150 28294 43218 28350
rect 43274 28294 43342 28350
rect 43398 28294 43494 28350
rect 42874 28226 43494 28294
rect 42874 28170 42970 28226
rect 43026 28170 43094 28226
rect 43150 28170 43218 28226
rect 43274 28170 43342 28226
rect 43398 28170 43494 28226
rect 42874 28102 43494 28170
rect 42874 28046 42970 28102
rect 43026 28046 43094 28102
rect 43150 28046 43218 28102
rect 43274 28046 43342 28102
rect 43398 28046 43494 28102
rect 42874 27978 43494 28046
rect 42874 27922 42970 27978
rect 43026 27922 43094 27978
rect 43150 27922 43218 27978
rect 43274 27922 43342 27978
rect 43398 27922 43494 27978
rect 42874 10350 43494 27922
rect 42874 10294 42970 10350
rect 43026 10294 43094 10350
rect 43150 10294 43218 10350
rect 43274 10294 43342 10350
rect 43398 10294 43494 10350
rect 42874 10226 43494 10294
rect 42874 10170 42970 10226
rect 43026 10170 43094 10226
rect 43150 10170 43218 10226
rect 43274 10170 43342 10226
rect 43398 10170 43494 10226
rect 42874 10102 43494 10170
rect 42874 10046 42970 10102
rect 43026 10046 43094 10102
rect 43150 10046 43218 10102
rect 43274 10046 43342 10102
rect 43398 10046 43494 10102
rect 42874 9978 43494 10046
rect 42874 9922 42970 9978
rect 43026 9922 43094 9978
rect 43150 9922 43218 9978
rect 43274 9922 43342 9978
rect 43398 9922 43494 9978
rect 42874 -1120 43494 9922
rect 42874 -1176 42970 -1120
rect 43026 -1176 43094 -1120
rect 43150 -1176 43218 -1120
rect 43274 -1176 43342 -1120
rect 43398 -1176 43494 -1120
rect 42874 -1244 43494 -1176
rect 42874 -1300 42970 -1244
rect 43026 -1300 43094 -1244
rect 43150 -1300 43218 -1244
rect 43274 -1300 43342 -1244
rect 43398 -1300 43494 -1244
rect 42874 -1368 43494 -1300
rect 42874 -1424 42970 -1368
rect 43026 -1424 43094 -1368
rect 43150 -1424 43218 -1368
rect 43274 -1424 43342 -1368
rect 43398 -1424 43494 -1368
rect 42874 -1492 43494 -1424
rect 42874 -1548 42970 -1492
rect 43026 -1548 43094 -1492
rect 43150 -1548 43218 -1492
rect 43274 -1548 43342 -1492
rect 43398 -1548 43494 -1492
rect 42874 -1644 43494 -1548
rect 57154 22350 57774 39922
rect 57154 22294 57250 22350
rect 57306 22294 57374 22350
rect 57430 22294 57498 22350
rect 57554 22294 57622 22350
rect 57678 22294 57774 22350
rect 57154 22226 57774 22294
rect 57154 22170 57250 22226
rect 57306 22170 57374 22226
rect 57430 22170 57498 22226
rect 57554 22170 57622 22226
rect 57678 22170 57774 22226
rect 57154 22102 57774 22170
rect 57154 22046 57250 22102
rect 57306 22046 57374 22102
rect 57430 22046 57498 22102
rect 57554 22046 57622 22102
rect 57678 22046 57774 22102
rect 57154 21978 57774 22046
rect 57154 21922 57250 21978
rect 57306 21922 57374 21978
rect 57430 21922 57498 21978
rect 57554 21922 57622 21978
rect 57678 21922 57774 21978
rect 57154 4350 57774 21922
rect 57154 4294 57250 4350
rect 57306 4294 57374 4350
rect 57430 4294 57498 4350
rect 57554 4294 57622 4350
rect 57678 4294 57774 4350
rect 57154 4226 57774 4294
rect 57154 4170 57250 4226
rect 57306 4170 57374 4226
rect 57430 4170 57498 4226
rect 57554 4170 57622 4226
rect 57678 4170 57774 4226
rect 57154 4102 57774 4170
rect 57154 4046 57250 4102
rect 57306 4046 57374 4102
rect 57430 4046 57498 4102
rect 57554 4046 57622 4102
rect 57678 4046 57774 4102
rect 57154 3978 57774 4046
rect 57154 3922 57250 3978
rect 57306 3922 57374 3978
rect 57430 3922 57498 3978
rect 57554 3922 57622 3978
rect 57678 3922 57774 3978
rect 57154 -160 57774 3922
rect 57154 -216 57250 -160
rect 57306 -216 57374 -160
rect 57430 -216 57498 -160
rect 57554 -216 57622 -160
rect 57678 -216 57774 -160
rect 57154 -284 57774 -216
rect 57154 -340 57250 -284
rect 57306 -340 57374 -284
rect 57430 -340 57498 -284
rect 57554 -340 57622 -284
rect 57678 -340 57774 -284
rect 57154 -408 57774 -340
rect 57154 -464 57250 -408
rect 57306 -464 57374 -408
rect 57430 -464 57498 -408
rect 57554 -464 57622 -408
rect 57678 -464 57774 -408
rect 57154 -532 57774 -464
rect 57154 -588 57250 -532
rect 57306 -588 57374 -532
rect 57430 -588 57498 -532
rect 57554 -588 57622 -532
rect 57678 -588 57774 -532
rect 57154 -1644 57774 -588
rect 60874 598172 61494 598268
rect 60874 598116 60970 598172
rect 61026 598116 61094 598172
rect 61150 598116 61218 598172
rect 61274 598116 61342 598172
rect 61398 598116 61494 598172
rect 60874 598048 61494 598116
rect 60874 597992 60970 598048
rect 61026 597992 61094 598048
rect 61150 597992 61218 598048
rect 61274 597992 61342 598048
rect 61398 597992 61494 598048
rect 60874 597924 61494 597992
rect 60874 597868 60970 597924
rect 61026 597868 61094 597924
rect 61150 597868 61218 597924
rect 61274 597868 61342 597924
rect 61398 597868 61494 597924
rect 60874 597800 61494 597868
rect 60874 597744 60970 597800
rect 61026 597744 61094 597800
rect 61150 597744 61218 597800
rect 61274 597744 61342 597800
rect 61398 597744 61494 597800
rect 60874 586350 61494 597744
rect 60874 586294 60970 586350
rect 61026 586294 61094 586350
rect 61150 586294 61218 586350
rect 61274 586294 61342 586350
rect 61398 586294 61494 586350
rect 60874 586226 61494 586294
rect 60874 586170 60970 586226
rect 61026 586170 61094 586226
rect 61150 586170 61218 586226
rect 61274 586170 61342 586226
rect 61398 586170 61494 586226
rect 60874 586102 61494 586170
rect 60874 586046 60970 586102
rect 61026 586046 61094 586102
rect 61150 586046 61218 586102
rect 61274 586046 61342 586102
rect 61398 586046 61494 586102
rect 60874 585978 61494 586046
rect 60874 585922 60970 585978
rect 61026 585922 61094 585978
rect 61150 585922 61218 585978
rect 61274 585922 61342 585978
rect 61398 585922 61494 585978
rect 60874 568350 61494 585922
rect 60874 568294 60970 568350
rect 61026 568294 61094 568350
rect 61150 568294 61218 568350
rect 61274 568294 61342 568350
rect 61398 568294 61494 568350
rect 60874 568226 61494 568294
rect 60874 568170 60970 568226
rect 61026 568170 61094 568226
rect 61150 568170 61218 568226
rect 61274 568170 61342 568226
rect 61398 568170 61494 568226
rect 60874 568102 61494 568170
rect 60874 568046 60970 568102
rect 61026 568046 61094 568102
rect 61150 568046 61218 568102
rect 61274 568046 61342 568102
rect 61398 568046 61494 568102
rect 60874 567978 61494 568046
rect 60874 567922 60970 567978
rect 61026 567922 61094 567978
rect 61150 567922 61218 567978
rect 61274 567922 61342 567978
rect 61398 567922 61494 567978
rect 60874 550350 61494 567922
rect 60874 550294 60970 550350
rect 61026 550294 61094 550350
rect 61150 550294 61218 550350
rect 61274 550294 61342 550350
rect 61398 550294 61494 550350
rect 60874 550226 61494 550294
rect 60874 550170 60970 550226
rect 61026 550170 61094 550226
rect 61150 550170 61218 550226
rect 61274 550170 61342 550226
rect 61398 550170 61494 550226
rect 60874 550102 61494 550170
rect 60874 550046 60970 550102
rect 61026 550046 61094 550102
rect 61150 550046 61218 550102
rect 61274 550046 61342 550102
rect 61398 550046 61494 550102
rect 60874 549978 61494 550046
rect 60874 549922 60970 549978
rect 61026 549922 61094 549978
rect 61150 549922 61218 549978
rect 61274 549922 61342 549978
rect 61398 549922 61494 549978
rect 60874 532350 61494 549922
rect 60874 532294 60970 532350
rect 61026 532294 61094 532350
rect 61150 532294 61218 532350
rect 61274 532294 61342 532350
rect 61398 532294 61494 532350
rect 60874 532226 61494 532294
rect 60874 532170 60970 532226
rect 61026 532170 61094 532226
rect 61150 532170 61218 532226
rect 61274 532170 61342 532226
rect 61398 532170 61494 532226
rect 60874 532102 61494 532170
rect 60874 532046 60970 532102
rect 61026 532046 61094 532102
rect 61150 532046 61218 532102
rect 61274 532046 61342 532102
rect 61398 532046 61494 532102
rect 60874 531978 61494 532046
rect 60874 531922 60970 531978
rect 61026 531922 61094 531978
rect 61150 531922 61218 531978
rect 61274 531922 61342 531978
rect 61398 531922 61494 531978
rect 60874 514350 61494 531922
rect 75154 597212 75774 598268
rect 75154 597156 75250 597212
rect 75306 597156 75374 597212
rect 75430 597156 75498 597212
rect 75554 597156 75622 597212
rect 75678 597156 75774 597212
rect 75154 597088 75774 597156
rect 75154 597032 75250 597088
rect 75306 597032 75374 597088
rect 75430 597032 75498 597088
rect 75554 597032 75622 597088
rect 75678 597032 75774 597088
rect 75154 596964 75774 597032
rect 75154 596908 75250 596964
rect 75306 596908 75374 596964
rect 75430 596908 75498 596964
rect 75554 596908 75622 596964
rect 75678 596908 75774 596964
rect 75154 596840 75774 596908
rect 75154 596784 75250 596840
rect 75306 596784 75374 596840
rect 75430 596784 75498 596840
rect 75554 596784 75622 596840
rect 75678 596784 75774 596840
rect 75154 580350 75774 596784
rect 75154 580294 75250 580350
rect 75306 580294 75374 580350
rect 75430 580294 75498 580350
rect 75554 580294 75622 580350
rect 75678 580294 75774 580350
rect 75154 580226 75774 580294
rect 75154 580170 75250 580226
rect 75306 580170 75374 580226
rect 75430 580170 75498 580226
rect 75554 580170 75622 580226
rect 75678 580170 75774 580226
rect 75154 580102 75774 580170
rect 75154 580046 75250 580102
rect 75306 580046 75374 580102
rect 75430 580046 75498 580102
rect 75554 580046 75622 580102
rect 75678 580046 75774 580102
rect 75154 579978 75774 580046
rect 75154 579922 75250 579978
rect 75306 579922 75374 579978
rect 75430 579922 75498 579978
rect 75554 579922 75622 579978
rect 75678 579922 75774 579978
rect 75154 562350 75774 579922
rect 75154 562294 75250 562350
rect 75306 562294 75374 562350
rect 75430 562294 75498 562350
rect 75554 562294 75622 562350
rect 75678 562294 75774 562350
rect 75154 562226 75774 562294
rect 75154 562170 75250 562226
rect 75306 562170 75374 562226
rect 75430 562170 75498 562226
rect 75554 562170 75622 562226
rect 75678 562170 75774 562226
rect 75154 562102 75774 562170
rect 75154 562046 75250 562102
rect 75306 562046 75374 562102
rect 75430 562046 75498 562102
rect 75554 562046 75622 562102
rect 75678 562046 75774 562102
rect 75154 561978 75774 562046
rect 75154 561922 75250 561978
rect 75306 561922 75374 561978
rect 75430 561922 75498 561978
rect 75554 561922 75622 561978
rect 75678 561922 75774 561978
rect 75154 544350 75774 561922
rect 75154 544294 75250 544350
rect 75306 544294 75374 544350
rect 75430 544294 75498 544350
rect 75554 544294 75622 544350
rect 75678 544294 75774 544350
rect 75154 544226 75774 544294
rect 75154 544170 75250 544226
rect 75306 544170 75374 544226
rect 75430 544170 75498 544226
rect 75554 544170 75622 544226
rect 75678 544170 75774 544226
rect 75154 544102 75774 544170
rect 75154 544046 75250 544102
rect 75306 544046 75374 544102
rect 75430 544046 75498 544102
rect 75554 544046 75622 544102
rect 75678 544046 75774 544102
rect 75154 543978 75774 544046
rect 75154 543922 75250 543978
rect 75306 543922 75374 543978
rect 75430 543922 75498 543978
rect 75554 543922 75622 543978
rect 75678 543922 75774 543978
rect 75154 526350 75774 543922
rect 75154 526294 75250 526350
rect 75306 526294 75374 526350
rect 75430 526294 75498 526350
rect 75554 526294 75622 526350
rect 75678 526294 75774 526350
rect 75154 526226 75774 526294
rect 75154 526170 75250 526226
rect 75306 526170 75374 526226
rect 75430 526170 75498 526226
rect 75554 526170 75622 526226
rect 75678 526170 75774 526226
rect 75154 526102 75774 526170
rect 75154 526046 75250 526102
rect 75306 526046 75374 526102
rect 75430 526046 75498 526102
rect 75554 526046 75622 526102
rect 75678 526046 75774 526102
rect 75154 525978 75774 526046
rect 75154 525922 75250 525978
rect 75306 525922 75374 525978
rect 75430 525922 75498 525978
rect 75554 525922 75622 525978
rect 75678 525922 75774 525978
rect 60874 514294 60970 514350
rect 61026 514294 61094 514350
rect 61150 514294 61218 514350
rect 61274 514294 61342 514350
rect 61398 514294 61494 514350
rect 60874 514226 61494 514294
rect 60874 514170 60970 514226
rect 61026 514170 61094 514226
rect 61150 514170 61218 514226
rect 61274 514170 61342 514226
rect 61398 514170 61494 514226
rect 60874 514102 61494 514170
rect 60874 514046 60970 514102
rect 61026 514046 61094 514102
rect 61150 514046 61218 514102
rect 61274 514046 61342 514102
rect 61398 514046 61494 514102
rect 60874 513978 61494 514046
rect 60874 513922 60970 513978
rect 61026 513922 61094 513978
rect 61150 513922 61218 513978
rect 61274 513922 61342 513978
rect 61398 513922 61494 513978
rect 60874 496350 61494 513922
rect 69808 514350 70128 514384
rect 69808 514294 69878 514350
rect 69934 514294 70002 514350
rect 70058 514294 70128 514350
rect 69808 514226 70128 514294
rect 69808 514170 69878 514226
rect 69934 514170 70002 514226
rect 70058 514170 70128 514226
rect 69808 514102 70128 514170
rect 69808 514046 69878 514102
rect 69934 514046 70002 514102
rect 70058 514046 70128 514102
rect 69808 513978 70128 514046
rect 69808 513922 69878 513978
rect 69934 513922 70002 513978
rect 70058 513922 70128 513978
rect 69808 513888 70128 513922
rect 75154 508350 75774 525922
rect 75154 508294 75250 508350
rect 75306 508294 75374 508350
rect 75430 508294 75498 508350
rect 75554 508294 75622 508350
rect 75678 508294 75774 508350
rect 75154 508226 75774 508294
rect 75154 508170 75250 508226
rect 75306 508170 75374 508226
rect 75430 508170 75498 508226
rect 75554 508170 75622 508226
rect 75678 508170 75774 508226
rect 75154 508102 75774 508170
rect 75154 508046 75250 508102
rect 75306 508046 75374 508102
rect 75430 508046 75498 508102
rect 75554 508046 75622 508102
rect 75678 508046 75774 508102
rect 75154 507978 75774 508046
rect 75154 507922 75250 507978
rect 75306 507922 75374 507978
rect 75430 507922 75498 507978
rect 75554 507922 75622 507978
rect 75678 507922 75774 507978
rect 60874 496294 60970 496350
rect 61026 496294 61094 496350
rect 61150 496294 61218 496350
rect 61274 496294 61342 496350
rect 61398 496294 61494 496350
rect 60874 496226 61494 496294
rect 60874 496170 60970 496226
rect 61026 496170 61094 496226
rect 61150 496170 61218 496226
rect 61274 496170 61342 496226
rect 61398 496170 61494 496226
rect 60874 496102 61494 496170
rect 60874 496046 60970 496102
rect 61026 496046 61094 496102
rect 61150 496046 61218 496102
rect 61274 496046 61342 496102
rect 61398 496046 61494 496102
rect 60874 495978 61494 496046
rect 60874 495922 60970 495978
rect 61026 495922 61094 495978
rect 61150 495922 61218 495978
rect 61274 495922 61342 495978
rect 61398 495922 61494 495978
rect 60874 478350 61494 495922
rect 69808 496350 70128 496384
rect 69808 496294 69878 496350
rect 69934 496294 70002 496350
rect 70058 496294 70128 496350
rect 69808 496226 70128 496294
rect 69808 496170 69878 496226
rect 69934 496170 70002 496226
rect 70058 496170 70128 496226
rect 69808 496102 70128 496170
rect 69808 496046 69878 496102
rect 69934 496046 70002 496102
rect 70058 496046 70128 496102
rect 69808 495978 70128 496046
rect 69808 495922 69878 495978
rect 69934 495922 70002 495978
rect 70058 495922 70128 495978
rect 69808 495888 70128 495922
rect 75154 490350 75774 507922
rect 75154 490294 75250 490350
rect 75306 490294 75374 490350
rect 75430 490294 75498 490350
rect 75554 490294 75622 490350
rect 75678 490294 75774 490350
rect 75154 490226 75774 490294
rect 75154 490170 75250 490226
rect 75306 490170 75374 490226
rect 75430 490170 75498 490226
rect 75554 490170 75622 490226
rect 75678 490170 75774 490226
rect 75154 490102 75774 490170
rect 75154 490046 75250 490102
rect 75306 490046 75374 490102
rect 75430 490046 75498 490102
rect 75554 490046 75622 490102
rect 75678 490046 75774 490102
rect 75154 489978 75774 490046
rect 75154 489922 75250 489978
rect 75306 489922 75374 489978
rect 75430 489922 75498 489978
rect 75554 489922 75622 489978
rect 75678 489922 75774 489978
rect 60874 478294 60970 478350
rect 61026 478294 61094 478350
rect 61150 478294 61218 478350
rect 61274 478294 61342 478350
rect 61398 478294 61494 478350
rect 60874 478226 61494 478294
rect 60874 478170 60970 478226
rect 61026 478170 61094 478226
rect 61150 478170 61218 478226
rect 61274 478170 61342 478226
rect 61398 478170 61494 478226
rect 60874 478102 61494 478170
rect 60874 478046 60970 478102
rect 61026 478046 61094 478102
rect 61150 478046 61218 478102
rect 61274 478046 61342 478102
rect 61398 478046 61494 478102
rect 60874 477978 61494 478046
rect 60874 477922 60970 477978
rect 61026 477922 61094 477978
rect 61150 477922 61218 477978
rect 61274 477922 61342 477978
rect 61398 477922 61494 477978
rect 60874 460350 61494 477922
rect 69808 478350 70128 478384
rect 69808 478294 69878 478350
rect 69934 478294 70002 478350
rect 70058 478294 70128 478350
rect 69808 478226 70128 478294
rect 69808 478170 69878 478226
rect 69934 478170 70002 478226
rect 70058 478170 70128 478226
rect 69808 478102 70128 478170
rect 69808 478046 69878 478102
rect 69934 478046 70002 478102
rect 70058 478046 70128 478102
rect 69808 477978 70128 478046
rect 69808 477922 69878 477978
rect 69934 477922 70002 477978
rect 70058 477922 70128 477978
rect 69808 477888 70128 477922
rect 75154 472350 75774 489922
rect 75154 472294 75250 472350
rect 75306 472294 75374 472350
rect 75430 472294 75498 472350
rect 75554 472294 75622 472350
rect 75678 472294 75774 472350
rect 75154 472226 75774 472294
rect 75154 472170 75250 472226
rect 75306 472170 75374 472226
rect 75430 472170 75498 472226
rect 75554 472170 75622 472226
rect 75678 472170 75774 472226
rect 75154 472102 75774 472170
rect 75154 472046 75250 472102
rect 75306 472046 75374 472102
rect 75430 472046 75498 472102
rect 75554 472046 75622 472102
rect 75678 472046 75774 472102
rect 75154 471978 75774 472046
rect 75154 471922 75250 471978
rect 75306 471922 75374 471978
rect 75430 471922 75498 471978
rect 75554 471922 75622 471978
rect 75678 471922 75774 471978
rect 60874 460294 60970 460350
rect 61026 460294 61094 460350
rect 61150 460294 61218 460350
rect 61274 460294 61342 460350
rect 61398 460294 61494 460350
rect 60874 460226 61494 460294
rect 60874 460170 60970 460226
rect 61026 460170 61094 460226
rect 61150 460170 61218 460226
rect 61274 460170 61342 460226
rect 61398 460170 61494 460226
rect 60874 460102 61494 460170
rect 60874 460046 60970 460102
rect 61026 460046 61094 460102
rect 61150 460046 61218 460102
rect 61274 460046 61342 460102
rect 61398 460046 61494 460102
rect 60874 459978 61494 460046
rect 60874 459922 60970 459978
rect 61026 459922 61094 459978
rect 61150 459922 61218 459978
rect 61274 459922 61342 459978
rect 61398 459922 61494 459978
rect 60874 442350 61494 459922
rect 69808 460350 70128 460384
rect 69808 460294 69878 460350
rect 69934 460294 70002 460350
rect 70058 460294 70128 460350
rect 69808 460226 70128 460294
rect 69808 460170 69878 460226
rect 69934 460170 70002 460226
rect 70058 460170 70128 460226
rect 69808 460102 70128 460170
rect 69808 460046 69878 460102
rect 69934 460046 70002 460102
rect 70058 460046 70128 460102
rect 69808 459978 70128 460046
rect 69808 459922 69878 459978
rect 69934 459922 70002 459978
rect 70058 459922 70128 459978
rect 69808 459888 70128 459922
rect 75154 454350 75774 471922
rect 75154 454294 75250 454350
rect 75306 454294 75374 454350
rect 75430 454294 75498 454350
rect 75554 454294 75622 454350
rect 75678 454294 75774 454350
rect 75154 454226 75774 454294
rect 75154 454170 75250 454226
rect 75306 454170 75374 454226
rect 75430 454170 75498 454226
rect 75554 454170 75622 454226
rect 75678 454170 75774 454226
rect 75154 454102 75774 454170
rect 75154 454046 75250 454102
rect 75306 454046 75374 454102
rect 75430 454046 75498 454102
rect 75554 454046 75622 454102
rect 75678 454046 75774 454102
rect 75154 453978 75774 454046
rect 75154 453922 75250 453978
rect 75306 453922 75374 453978
rect 75430 453922 75498 453978
rect 75554 453922 75622 453978
rect 75678 453922 75774 453978
rect 60874 442294 60970 442350
rect 61026 442294 61094 442350
rect 61150 442294 61218 442350
rect 61274 442294 61342 442350
rect 61398 442294 61494 442350
rect 60874 442226 61494 442294
rect 60874 442170 60970 442226
rect 61026 442170 61094 442226
rect 61150 442170 61218 442226
rect 61274 442170 61342 442226
rect 61398 442170 61494 442226
rect 60874 442102 61494 442170
rect 60874 442046 60970 442102
rect 61026 442046 61094 442102
rect 61150 442046 61218 442102
rect 61274 442046 61342 442102
rect 61398 442046 61494 442102
rect 60874 441978 61494 442046
rect 60874 441922 60970 441978
rect 61026 441922 61094 441978
rect 61150 441922 61218 441978
rect 61274 441922 61342 441978
rect 61398 441922 61494 441978
rect 60874 424350 61494 441922
rect 69808 442350 70128 442384
rect 69808 442294 69878 442350
rect 69934 442294 70002 442350
rect 70058 442294 70128 442350
rect 69808 442226 70128 442294
rect 69808 442170 69878 442226
rect 69934 442170 70002 442226
rect 70058 442170 70128 442226
rect 69808 442102 70128 442170
rect 69808 442046 69878 442102
rect 69934 442046 70002 442102
rect 70058 442046 70128 442102
rect 69808 441978 70128 442046
rect 69808 441922 69878 441978
rect 69934 441922 70002 441978
rect 70058 441922 70128 441978
rect 69808 441888 70128 441922
rect 75154 436350 75774 453922
rect 75154 436294 75250 436350
rect 75306 436294 75374 436350
rect 75430 436294 75498 436350
rect 75554 436294 75622 436350
rect 75678 436294 75774 436350
rect 75154 436226 75774 436294
rect 75154 436170 75250 436226
rect 75306 436170 75374 436226
rect 75430 436170 75498 436226
rect 75554 436170 75622 436226
rect 75678 436170 75774 436226
rect 75154 436102 75774 436170
rect 75154 436046 75250 436102
rect 75306 436046 75374 436102
rect 75430 436046 75498 436102
rect 75554 436046 75622 436102
rect 75678 436046 75774 436102
rect 75154 435978 75774 436046
rect 75154 435922 75250 435978
rect 75306 435922 75374 435978
rect 75430 435922 75498 435978
rect 75554 435922 75622 435978
rect 75678 435922 75774 435978
rect 60874 424294 60970 424350
rect 61026 424294 61094 424350
rect 61150 424294 61218 424350
rect 61274 424294 61342 424350
rect 61398 424294 61494 424350
rect 60874 424226 61494 424294
rect 60874 424170 60970 424226
rect 61026 424170 61094 424226
rect 61150 424170 61218 424226
rect 61274 424170 61342 424226
rect 61398 424170 61494 424226
rect 60874 424102 61494 424170
rect 60874 424046 60970 424102
rect 61026 424046 61094 424102
rect 61150 424046 61218 424102
rect 61274 424046 61342 424102
rect 61398 424046 61494 424102
rect 60874 423978 61494 424046
rect 60874 423922 60970 423978
rect 61026 423922 61094 423978
rect 61150 423922 61218 423978
rect 61274 423922 61342 423978
rect 61398 423922 61494 423978
rect 60874 406350 61494 423922
rect 69808 424350 70128 424384
rect 69808 424294 69878 424350
rect 69934 424294 70002 424350
rect 70058 424294 70128 424350
rect 69808 424226 70128 424294
rect 69808 424170 69878 424226
rect 69934 424170 70002 424226
rect 70058 424170 70128 424226
rect 69808 424102 70128 424170
rect 69808 424046 69878 424102
rect 69934 424046 70002 424102
rect 70058 424046 70128 424102
rect 69808 423978 70128 424046
rect 69808 423922 69878 423978
rect 69934 423922 70002 423978
rect 70058 423922 70128 423978
rect 69808 423888 70128 423922
rect 75154 418350 75774 435922
rect 75154 418294 75250 418350
rect 75306 418294 75374 418350
rect 75430 418294 75498 418350
rect 75554 418294 75622 418350
rect 75678 418294 75774 418350
rect 75154 418226 75774 418294
rect 75154 418170 75250 418226
rect 75306 418170 75374 418226
rect 75430 418170 75498 418226
rect 75554 418170 75622 418226
rect 75678 418170 75774 418226
rect 75154 418102 75774 418170
rect 75154 418046 75250 418102
rect 75306 418046 75374 418102
rect 75430 418046 75498 418102
rect 75554 418046 75622 418102
rect 75678 418046 75774 418102
rect 75154 417978 75774 418046
rect 75154 417922 75250 417978
rect 75306 417922 75374 417978
rect 75430 417922 75498 417978
rect 75554 417922 75622 417978
rect 75678 417922 75774 417978
rect 60874 406294 60970 406350
rect 61026 406294 61094 406350
rect 61150 406294 61218 406350
rect 61274 406294 61342 406350
rect 61398 406294 61494 406350
rect 60874 406226 61494 406294
rect 60874 406170 60970 406226
rect 61026 406170 61094 406226
rect 61150 406170 61218 406226
rect 61274 406170 61342 406226
rect 61398 406170 61494 406226
rect 60874 406102 61494 406170
rect 60874 406046 60970 406102
rect 61026 406046 61094 406102
rect 61150 406046 61218 406102
rect 61274 406046 61342 406102
rect 61398 406046 61494 406102
rect 60874 405978 61494 406046
rect 60874 405922 60970 405978
rect 61026 405922 61094 405978
rect 61150 405922 61218 405978
rect 61274 405922 61342 405978
rect 61398 405922 61494 405978
rect 60874 388350 61494 405922
rect 69808 406350 70128 406384
rect 69808 406294 69878 406350
rect 69934 406294 70002 406350
rect 70058 406294 70128 406350
rect 69808 406226 70128 406294
rect 69808 406170 69878 406226
rect 69934 406170 70002 406226
rect 70058 406170 70128 406226
rect 69808 406102 70128 406170
rect 69808 406046 69878 406102
rect 69934 406046 70002 406102
rect 70058 406046 70128 406102
rect 69808 405978 70128 406046
rect 69808 405922 69878 405978
rect 69934 405922 70002 405978
rect 70058 405922 70128 405978
rect 69808 405888 70128 405922
rect 75154 400350 75774 417922
rect 75154 400294 75250 400350
rect 75306 400294 75374 400350
rect 75430 400294 75498 400350
rect 75554 400294 75622 400350
rect 75678 400294 75774 400350
rect 75154 400226 75774 400294
rect 75154 400170 75250 400226
rect 75306 400170 75374 400226
rect 75430 400170 75498 400226
rect 75554 400170 75622 400226
rect 75678 400170 75774 400226
rect 75154 400102 75774 400170
rect 75154 400046 75250 400102
rect 75306 400046 75374 400102
rect 75430 400046 75498 400102
rect 75554 400046 75622 400102
rect 75678 400046 75774 400102
rect 75154 399978 75774 400046
rect 75154 399922 75250 399978
rect 75306 399922 75374 399978
rect 75430 399922 75498 399978
rect 75554 399922 75622 399978
rect 75678 399922 75774 399978
rect 60874 388294 60970 388350
rect 61026 388294 61094 388350
rect 61150 388294 61218 388350
rect 61274 388294 61342 388350
rect 61398 388294 61494 388350
rect 60874 388226 61494 388294
rect 60874 388170 60970 388226
rect 61026 388170 61094 388226
rect 61150 388170 61218 388226
rect 61274 388170 61342 388226
rect 61398 388170 61494 388226
rect 60874 388102 61494 388170
rect 60874 388046 60970 388102
rect 61026 388046 61094 388102
rect 61150 388046 61218 388102
rect 61274 388046 61342 388102
rect 61398 388046 61494 388102
rect 60874 387978 61494 388046
rect 60874 387922 60970 387978
rect 61026 387922 61094 387978
rect 61150 387922 61218 387978
rect 61274 387922 61342 387978
rect 61398 387922 61494 387978
rect 60874 370350 61494 387922
rect 69808 388350 70128 388384
rect 69808 388294 69878 388350
rect 69934 388294 70002 388350
rect 70058 388294 70128 388350
rect 69808 388226 70128 388294
rect 69808 388170 69878 388226
rect 69934 388170 70002 388226
rect 70058 388170 70128 388226
rect 69808 388102 70128 388170
rect 69808 388046 69878 388102
rect 69934 388046 70002 388102
rect 70058 388046 70128 388102
rect 69808 387978 70128 388046
rect 69808 387922 69878 387978
rect 69934 387922 70002 387978
rect 70058 387922 70128 387978
rect 69808 387888 70128 387922
rect 75154 382350 75774 399922
rect 75154 382294 75250 382350
rect 75306 382294 75374 382350
rect 75430 382294 75498 382350
rect 75554 382294 75622 382350
rect 75678 382294 75774 382350
rect 75154 382226 75774 382294
rect 75154 382170 75250 382226
rect 75306 382170 75374 382226
rect 75430 382170 75498 382226
rect 75554 382170 75622 382226
rect 75678 382170 75774 382226
rect 75154 382102 75774 382170
rect 75154 382046 75250 382102
rect 75306 382046 75374 382102
rect 75430 382046 75498 382102
rect 75554 382046 75622 382102
rect 75678 382046 75774 382102
rect 75154 381978 75774 382046
rect 75154 381922 75250 381978
rect 75306 381922 75374 381978
rect 75430 381922 75498 381978
rect 75554 381922 75622 381978
rect 75678 381922 75774 381978
rect 60874 370294 60970 370350
rect 61026 370294 61094 370350
rect 61150 370294 61218 370350
rect 61274 370294 61342 370350
rect 61398 370294 61494 370350
rect 60874 370226 61494 370294
rect 60874 370170 60970 370226
rect 61026 370170 61094 370226
rect 61150 370170 61218 370226
rect 61274 370170 61342 370226
rect 61398 370170 61494 370226
rect 60874 370102 61494 370170
rect 60874 370046 60970 370102
rect 61026 370046 61094 370102
rect 61150 370046 61218 370102
rect 61274 370046 61342 370102
rect 61398 370046 61494 370102
rect 60874 369978 61494 370046
rect 60874 369922 60970 369978
rect 61026 369922 61094 369978
rect 61150 369922 61218 369978
rect 61274 369922 61342 369978
rect 61398 369922 61494 369978
rect 60874 352350 61494 369922
rect 69808 370350 70128 370384
rect 69808 370294 69878 370350
rect 69934 370294 70002 370350
rect 70058 370294 70128 370350
rect 69808 370226 70128 370294
rect 69808 370170 69878 370226
rect 69934 370170 70002 370226
rect 70058 370170 70128 370226
rect 69808 370102 70128 370170
rect 69808 370046 69878 370102
rect 69934 370046 70002 370102
rect 70058 370046 70128 370102
rect 69808 369978 70128 370046
rect 69808 369922 69878 369978
rect 69934 369922 70002 369978
rect 70058 369922 70128 369978
rect 69808 369888 70128 369922
rect 75154 364350 75774 381922
rect 75154 364294 75250 364350
rect 75306 364294 75374 364350
rect 75430 364294 75498 364350
rect 75554 364294 75622 364350
rect 75678 364294 75774 364350
rect 75154 364226 75774 364294
rect 75154 364170 75250 364226
rect 75306 364170 75374 364226
rect 75430 364170 75498 364226
rect 75554 364170 75622 364226
rect 75678 364170 75774 364226
rect 75154 364102 75774 364170
rect 75154 364046 75250 364102
rect 75306 364046 75374 364102
rect 75430 364046 75498 364102
rect 75554 364046 75622 364102
rect 75678 364046 75774 364102
rect 75154 363978 75774 364046
rect 75154 363922 75250 363978
rect 75306 363922 75374 363978
rect 75430 363922 75498 363978
rect 75554 363922 75622 363978
rect 75678 363922 75774 363978
rect 60874 352294 60970 352350
rect 61026 352294 61094 352350
rect 61150 352294 61218 352350
rect 61274 352294 61342 352350
rect 61398 352294 61494 352350
rect 60874 352226 61494 352294
rect 60874 352170 60970 352226
rect 61026 352170 61094 352226
rect 61150 352170 61218 352226
rect 61274 352170 61342 352226
rect 61398 352170 61494 352226
rect 60874 352102 61494 352170
rect 60874 352046 60970 352102
rect 61026 352046 61094 352102
rect 61150 352046 61218 352102
rect 61274 352046 61342 352102
rect 61398 352046 61494 352102
rect 60874 351978 61494 352046
rect 60874 351922 60970 351978
rect 61026 351922 61094 351978
rect 61150 351922 61218 351978
rect 61274 351922 61342 351978
rect 61398 351922 61494 351978
rect 60874 334350 61494 351922
rect 69808 352350 70128 352384
rect 69808 352294 69878 352350
rect 69934 352294 70002 352350
rect 70058 352294 70128 352350
rect 69808 352226 70128 352294
rect 69808 352170 69878 352226
rect 69934 352170 70002 352226
rect 70058 352170 70128 352226
rect 69808 352102 70128 352170
rect 69808 352046 69878 352102
rect 69934 352046 70002 352102
rect 70058 352046 70128 352102
rect 69808 351978 70128 352046
rect 69808 351922 69878 351978
rect 69934 351922 70002 351978
rect 70058 351922 70128 351978
rect 69808 351888 70128 351922
rect 75154 346350 75774 363922
rect 75154 346294 75250 346350
rect 75306 346294 75374 346350
rect 75430 346294 75498 346350
rect 75554 346294 75622 346350
rect 75678 346294 75774 346350
rect 75154 346226 75774 346294
rect 75154 346170 75250 346226
rect 75306 346170 75374 346226
rect 75430 346170 75498 346226
rect 75554 346170 75622 346226
rect 75678 346170 75774 346226
rect 75154 346102 75774 346170
rect 75154 346046 75250 346102
rect 75306 346046 75374 346102
rect 75430 346046 75498 346102
rect 75554 346046 75622 346102
rect 75678 346046 75774 346102
rect 75154 345978 75774 346046
rect 75154 345922 75250 345978
rect 75306 345922 75374 345978
rect 75430 345922 75498 345978
rect 75554 345922 75622 345978
rect 75678 345922 75774 345978
rect 60874 334294 60970 334350
rect 61026 334294 61094 334350
rect 61150 334294 61218 334350
rect 61274 334294 61342 334350
rect 61398 334294 61494 334350
rect 60874 334226 61494 334294
rect 60874 334170 60970 334226
rect 61026 334170 61094 334226
rect 61150 334170 61218 334226
rect 61274 334170 61342 334226
rect 61398 334170 61494 334226
rect 60874 334102 61494 334170
rect 60874 334046 60970 334102
rect 61026 334046 61094 334102
rect 61150 334046 61218 334102
rect 61274 334046 61342 334102
rect 61398 334046 61494 334102
rect 60874 333978 61494 334046
rect 60874 333922 60970 333978
rect 61026 333922 61094 333978
rect 61150 333922 61218 333978
rect 61274 333922 61342 333978
rect 61398 333922 61494 333978
rect 60874 316350 61494 333922
rect 69808 334350 70128 334384
rect 69808 334294 69878 334350
rect 69934 334294 70002 334350
rect 70058 334294 70128 334350
rect 69808 334226 70128 334294
rect 69808 334170 69878 334226
rect 69934 334170 70002 334226
rect 70058 334170 70128 334226
rect 69808 334102 70128 334170
rect 69808 334046 69878 334102
rect 69934 334046 70002 334102
rect 70058 334046 70128 334102
rect 69808 333978 70128 334046
rect 69808 333922 69878 333978
rect 69934 333922 70002 333978
rect 70058 333922 70128 333978
rect 69808 333888 70128 333922
rect 75154 328350 75774 345922
rect 75154 328294 75250 328350
rect 75306 328294 75374 328350
rect 75430 328294 75498 328350
rect 75554 328294 75622 328350
rect 75678 328294 75774 328350
rect 75154 328226 75774 328294
rect 75154 328170 75250 328226
rect 75306 328170 75374 328226
rect 75430 328170 75498 328226
rect 75554 328170 75622 328226
rect 75678 328170 75774 328226
rect 75154 328102 75774 328170
rect 75154 328046 75250 328102
rect 75306 328046 75374 328102
rect 75430 328046 75498 328102
rect 75554 328046 75622 328102
rect 75678 328046 75774 328102
rect 75154 327978 75774 328046
rect 75154 327922 75250 327978
rect 75306 327922 75374 327978
rect 75430 327922 75498 327978
rect 75554 327922 75622 327978
rect 75678 327922 75774 327978
rect 60874 316294 60970 316350
rect 61026 316294 61094 316350
rect 61150 316294 61218 316350
rect 61274 316294 61342 316350
rect 61398 316294 61494 316350
rect 60874 316226 61494 316294
rect 60874 316170 60970 316226
rect 61026 316170 61094 316226
rect 61150 316170 61218 316226
rect 61274 316170 61342 316226
rect 61398 316170 61494 316226
rect 60874 316102 61494 316170
rect 60874 316046 60970 316102
rect 61026 316046 61094 316102
rect 61150 316046 61218 316102
rect 61274 316046 61342 316102
rect 61398 316046 61494 316102
rect 60874 315978 61494 316046
rect 60874 315922 60970 315978
rect 61026 315922 61094 315978
rect 61150 315922 61218 315978
rect 61274 315922 61342 315978
rect 61398 315922 61494 315978
rect 60874 298350 61494 315922
rect 69808 316350 70128 316384
rect 69808 316294 69878 316350
rect 69934 316294 70002 316350
rect 70058 316294 70128 316350
rect 69808 316226 70128 316294
rect 69808 316170 69878 316226
rect 69934 316170 70002 316226
rect 70058 316170 70128 316226
rect 69808 316102 70128 316170
rect 69808 316046 69878 316102
rect 69934 316046 70002 316102
rect 70058 316046 70128 316102
rect 69808 315978 70128 316046
rect 69808 315922 69878 315978
rect 69934 315922 70002 315978
rect 70058 315922 70128 315978
rect 69808 315888 70128 315922
rect 75154 310350 75774 327922
rect 75154 310294 75250 310350
rect 75306 310294 75374 310350
rect 75430 310294 75498 310350
rect 75554 310294 75622 310350
rect 75678 310294 75774 310350
rect 75154 310226 75774 310294
rect 75154 310170 75250 310226
rect 75306 310170 75374 310226
rect 75430 310170 75498 310226
rect 75554 310170 75622 310226
rect 75678 310170 75774 310226
rect 75154 310102 75774 310170
rect 75154 310046 75250 310102
rect 75306 310046 75374 310102
rect 75430 310046 75498 310102
rect 75554 310046 75622 310102
rect 75678 310046 75774 310102
rect 75154 309978 75774 310046
rect 75154 309922 75250 309978
rect 75306 309922 75374 309978
rect 75430 309922 75498 309978
rect 75554 309922 75622 309978
rect 75678 309922 75774 309978
rect 60874 298294 60970 298350
rect 61026 298294 61094 298350
rect 61150 298294 61218 298350
rect 61274 298294 61342 298350
rect 61398 298294 61494 298350
rect 60874 298226 61494 298294
rect 60874 298170 60970 298226
rect 61026 298170 61094 298226
rect 61150 298170 61218 298226
rect 61274 298170 61342 298226
rect 61398 298170 61494 298226
rect 60874 298102 61494 298170
rect 60874 298046 60970 298102
rect 61026 298046 61094 298102
rect 61150 298046 61218 298102
rect 61274 298046 61342 298102
rect 61398 298046 61494 298102
rect 60874 297978 61494 298046
rect 60874 297922 60970 297978
rect 61026 297922 61094 297978
rect 61150 297922 61218 297978
rect 61274 297922 61342 297978
rect 61398 297922 61494 297978
rect 60874 280350 61494 297922
rect 69808 298350 70128 298384
rect 69808 298294 69878 298350
rect 69934 298294 70002 298350
rect 70058 298294 70128 298350
rect 69808 298226 70128 298294
rect 69808 298170 69878 298226
rect 69934 298170 70002 298226
rect 70058 298170 70128 298226
rect 69808 298102 70128 298170
rect 69808 298046 69878 298102
rect 69934 298046 70002 298102
rect 70058 298046 70128 298102
rect 69808 297978 70128 298046
rect 69808 297922 69878 297978
rect 69934 297922 70002 297978
rect 70058 297922 70128 297978
rect 69808 297888 70128 297922
rect 75154 292350 75774 309922
rect 75154 292294 75250 292350
rect 75306 292294 75374 292350
rect 75430 292294 75498 292350
rect 75554 292294 75622 292350
rect 75678 292294 75774 292350
rect 75154 292226 75774 292294
rect 75154 292170 75250 292226
rect 75306 292170 75374 292226
rect 75430 292170 75498 292226
rect 75554 292170 75622 292226
rect 75678 292170 75774 292226
rect 75154 292102 75774 292170
rect 75154 292046 75250 292102
rect 75306 292046 75374 292102
rect 75430 292046 75498 292102
rect 75554 292046 75622 292102
rect 75678 292046 75774 292102
rect 75154 291978 75774 292046
rect 75154 291922 75250 291978
rect 75306 291922 75374 291978
rect 75430 291922 75498 291978
rect 75554 291922 75622 291978
rect 75678 291922 75774 291978
rect 60874 280294 60970 280350
rect 61026 280294 61094 280350
rect 61150 280294 61218 280350
rect 61274 280294 61342 280350
rect 61398 280294 61494 280350
rect 60874 280226 61494 280294
rect 60874 280170 60970 280226
rect 61026 280170 61094 280226
rect 61150 280170 61218 280226
rect 61274 280170 61342 280226
rect 61398 280170 61494 280226
rect 60874 280102 61494 280170
rect 60874 280046 60970 280102
rect 61026 280046 61094 280102
rect 61150 280046 61218 280102
rect 61274 280046 61342 280102
rect 61398 280046 61494 280102
rect 60874 279978 61494 280046
rect 60874 279922 60970 279978
rect 61026 279922 61094 279978
rect 61150 279922 61218 279978
rect 61274 279922 61342 279978
rect 61398 279922 61494 279978
rect 60874 262350 61494 279922
rect 69808 280350 70128 280384
rect 69808 280294 69878 280350
rect 69934 280294 70002 280350
rect 70058 280294 70128 280350
rect 69808 280226 70128 280294
rect 69808 280170 69878 280226
rect 69934 280170 70002 280226
rect 70058 280170 70128 280226
rect 69808 280102 70128 280170
rect 69808 280046 69878 280102
rect 69934 280046 70002 280102
rect 70058 280046 70128 280102
rect 69808 279978 70128 280046
rect 69808 279922 69878 279978
rect 69934 279922 70002 279978
rect 70058 279922 70128 279978
rect 69808 279888 70128 279922
rect 75154 274350 75774 291922
rect 75154 274294 75250 274350
rect 75306 274294 75374 274350
rect 75430 274294 75498 274350
rect 75554 274294 75622 274350
rect 75678 274294 75774 274350
rect 75154 274226 75774 274294
rect 75154 274170 75250 274226
rect 75306 274170 75374 274226
rect 75430 274170 75498 274226
rect 75554 274170 75622 274226
rect 75678 274170 75774 274226
rect 75154 274102 75774 274170
rect 75154 274046 75250 274102
rect 75306 274046 75374 274102
rect 75430 274046 75498 274102
rect 75554 274046 75622 274102
rect 75678 274046 75774 274102
rect 75154 273978 75774 274046
rect 75154 273922 75250 273978
rect 75306 273922 75374 273978
rect 75430 273922 75498 273978
rect 75554 273922 75622 273978
rect 75678 273922 75774 273978
rect 60874 262294 60970 262350
rect 61026 262294 61094 262350
rect 61150 262294 61218 262350
rect 61274 262294 61342 262350
rect 61398 262294 61494 262350
rect 60874 262226 61494 262294
rect 60874 262170 60970 262226
rect 61026 262170 61094 262226
rect 61150 262170 61218 262226
rect 61274 262170 61342 262226
rect 61398 262170 61494 262226
rect 60874 262102 61494 262170
rect 60874 262046 60970 262102
rect 61026 262046 61094 262102
rect 61150 262046 61218 262102
rect 61274 262046 61342 262102
rect 61398 262046 61494 262102
rect 60874 261978 61494 262046
rect 60874 261922 60970 261978
rect 61026 261922 61094 261978
rect 61150 261922 61218 261978
rect 61274 261922 61342 261978
rect 61398 261922 61494 261978
rect 60874 244350 61494 261922
rect 69808 262350 70128 262384
rect 69808 262294 69878 262350
rect 69934 262294 70002 262350
rect 70058 262294 70128 262350
rect 69808 262226 70128 262294
rect 69808 262170 69878 262226
rect 69934 262170 70002 262226
rect 70058 262170 70128 262226
rect 69808 262102 70128 262170
rect 69808 262046 69878 262102
rect 69934 262046 70002 262102
rect 70058 262046 70128 262102
rect 69808 261978 70128 262046
rect 69808 261922 69878 261978
rect 69934 261922 70002 261978
rect 70058 261922 70128 261978
rect 69808 261888 70128 261922
rect 75154 256350 75774 273922
rect 75154 256294 75250 256350
rect 75306 256294 75374 256350
rect 75430 256294 75498 256350
rect 75554 256294 75622 256350
rect 75678 256294 75774 256350
rect 75154 256226 75774 256294
rect 75154 256170 75250 256226
rect 75306 256170 75374 256226
rect 75430 256170 75498 256226
rect 75554 256170 75622 256226
rect 75678 256170 75774 256226
rect 75154 256102 75774 256170
rect 75154 256046 75250 256102
rect 75306 256046 75374 256102
rect 75430 256046 75498 256102
rect 75554 256046 75622 256102
rect 75678 256046 75774 256102
rect 75154 255978 75774 256046
rect 75154 255922 75250 255978
rect 75306 255922 75374 255978
rect 75430 255922 75498 255978
rect 75554 255922 75622 255978
rect 75678 255922 75774 255978
rect 60874 244294 60970 244350
rect 61026 244294 61094 244350
rect 61150 244294 61218 244350
rect 61274 244294 61342 244350
rect 61398 244294 61494 244350
rect 60874 244226 61494 244294
rect 60874 244170 60970 244226
rect 61026 244170 61094 244226
rect 61150 244170 61218 244226
rect 61274 244170 61342 244226
rect 61398 244170 61494 244226
rect 60874 244102 61494 244170
rect 60874 244046 60970 244102
rect 61026 244046 61094 244102
rect 61150 244046 61218 244102
rect 61274 244046 61342 244102
rect 61398 244046 61494 244102
rect 60874 243978 61494 244046
rect 60874 243922 60970 243978
rect 61026 243922 61094 243978
rect 61150 243922 61218 243978
rect 61274 243922 61342 243978
rect 61398 243922 61494 243978
rect 60874 226350 61494 243922
rect 69808 244350 70128 244384
rect 69808 244294 69878 244350
rect 69934 244294 70002 244350
rect 70058 244294 70128 244350
rect 69808 244226 70128 244294
rect 69808 244170 69878 244226
rect 69934 244170 70002 244226
rect 70058 244170 70128 244226
rect 69808 244102 70128 244170
rect 69808 244046 69878 244102
rect 69934 244046 70002 244102
rect 70058 244046 70128 244102
rect 69808 243978 70128 244046
rect 69808 243922 69878 243978
rect 69934 243922 70002 243978
rect 70058 243922 70128 243978
rect 69808 243888 70128 243922
rect 75154 238350 75774 255922
rect 75154 238294 75250 238350
rect 75306 238294 75374 238350
rect 75430 238294 75498 238350
rect 75554 238294 75622 238350
rect 75678 238294 75774 238350
rect 75154 238226 75774 238294
rect 75154 238170 75250 238226
rect 75306 238170 75374 238226
rect 75430 238170 75498 238226
rect 75554 238170 75622 238226
rect 75678 238170 75774 238226
rect 75154 238102 75774 238170
rect 75154 238046 75250 238102
rect 75306 238046 75374 238102
rect 75430 238046 75498 238102
rect 75554 238046 75622 238102
rect 75678 238046 75774 238102
rect 75154 237978 75774 238046
rect 75154 237922 75250 237978
rect 75306 237922 75374 237978
rect 75430 237922 75498 237978
rect 75554 237922 75622 237978
rect 75678 237922 75774 237978
rect 60874 226294 60970 226350
rect 61026 226294 61094 226350
rect 61150 226294 61218 226350
rect 61274 226294 61342 226350
rect 61398 226294 61494 226350
rect 60874 226226 61494 226294
rect 60874 226170 60970 226226
rect 61026 226170 61094 226226
rect 61150 226170 61218 226226
rect 61274 226170 61342 226226
rect 61398 226170 61494 226226
rect 60874 226102 61494 226170
rect 60874 226046 60970 226102
rect 61026 226046 61094 226102
rect 61150 226046 61218 226102
rect 61274 226046 61342 226102
rect 61398 226046 61494 226102
rect 60874 225978 61494 226046
rect 60874 225922 60970 225978
rect 61026 225922 61094 225978
rect 61150 225922 61218 225978
rect 61274 225922 61342 225978
rect 61398 225922 61494 225978
rect 60874 208350 61494 225922
rect 69808 226350 70128 226384
rect 69808 226294 69878 226350
rect 69934 226294 70002 226350
rect 70058 226294 70128 226350
rect 69808 226226 70128 226294
rect 69808 226170 69878 226226
rect 69934 226170 70002 226226
rect 70058 226170 70128 226226
rect 69808 226102 70128 226170
rect 69808 226046 69878 226102
rect 69934 226046 70002 226102
rect 70058 226046 70128 226102
rect 69808 225978 70128 226046
rect 69808 225922 69878 225978
rect 69934 225922 70002 225978
rect 70058 225922 70128 225978
rect 69808 225888 70128 225922
rect 75154 220350 75774 237922
rect 75154 220294 75250 220350
rect 75306 220294 75374 220350
rect 75430 220294 75498 220350
rect 75554 220294 75622 220350
rect 75678 220294 75774 220350
rect 75154 220226 75774 220294
rect 75154 220170 75250 220226
rect 75306 220170 75374 220226
rect 75430 220170 75498 220226
rect 75554 220170 75622 220226
rect 75678 220170 75774 220226
rect 75154 220102 75774 220170
rect 75154 220046 75250 220102
rect 75306 220046 75374 220102
rect 75430 220046 75498 220102
rect 75554 220046 75622 220102
rect 75678 220046 75774 220102
rect 75154 219978 75774 220046
rect 75154 219922 75250 219978
rect 75306 219922 75374 219978
rect 75430 219922 75498 219978
rect 75554 219922 75622 219978
rect 75678 219922 75774 219978
rect 60874 208294 60970 208350
rect 61026 208294 61094 208350
rect 61150 208294 61218 208350
rect 61274 208294 61342 208350
rect 61398 208294 61494 208350
rect 60874 208226 61494 208294
rect 60874 208170 60970 208226
rect 61026 208170 61094 208226
rect 61150 208170 61218 208226
rect 61274 208170 61342 208226
rect 61398 208170 61494 208226
rect 60874 208102 61494 208170
rect 60874 208046 60970 208102
rect 61026 208046 61094 208102
rect 61150 208046 61218 208102
rect 61274 208046 61342 208102
rect 61398 208046 61494 208102
rect 60874 207978 61494 208046
rect 60874 207922 60970 207978
rect 61026 207922 61094 207978
rect 61150 207922 61218 207978
rect 61274 207922 61342 207978
rect 61398 207922 61494 207978
rect 60874 190350 61494 207922
rect 69808 208350 70128 208384
rect 69808 208294 69878 208350
rect 69934 208294 70002 208350
rect 70058 208294 70128 208350
rect 69808 208226 70128 208294
rect 69808 208170 69878 208226
rect 69934 208170 70002 208226
rect 70058 208170 70128 208226
rect 69808 208102 70128 208170
rect 69808 208046 69878 208102
rect 69934 208046 70002 208102
rect 70058 208046 70128 208102
rect 69808 207978 70128 208046
rect 69808 207922 69878 207978
rect 69934 207922 70002 207978
rect 70058 207922 70128 207978
rect 69808 207888 70128 207922
rect 75154 202350 75774 219922
rect 75154 202294 75250 202350
rect 75306 202294 75374 202350
rect 75430 202294 75498 202350
rect 75554 202294 75622 202350
rect 75678 202294 75774 202350
rect 75154 202226 75774 202294
rect 75154 202170 75250 202226
rect 75306 202170 75374 202226
rect 75430 202170 75498 202226
rect 75554 202170 75622 202226
rect 75678 202170 75774 202226
rect 75154 202102 75774 202170
rect 75154 202046 75250 202102
rect 75306 202046 75374 202102
rect 75430 202046 75498 202102
rect 75554 202046 75622 202102
rect 75678 202046 75774 202102
rect 75154 201978 75774 202046
rect 75154 201922 75250 201978
rect 75306 201922 75374 201978
rect 75430 201922 75498 201978
rect 75554 201922 75622 201978
rect 75678 201922 75774 201978
rect 60874 190294 60970 190350
rect 61026 190294 61094 190350
rect 61150 190294 61218 190350
rect 61274 190294 61342 190350
rect 61398 190294 61494 190350
rect 60874 190226 61494 190294
rect 60874 190170 60970 190226
rect 61026 190170 61094 190226
rect 61150 190170 61218 190226
rect 61274 190170 61342 190226
rect 61398 190170 61494 190226
rect 60874 190102 61494 190170
rect 60874 190046 60970 190102
rect 61026 190046 61094 190102
rect 61150 190046 61218 190102
rect 61274 190046 61342 190102
rect 61398 190046 61494 190102
rect 60874 189978 61494 190046
rect 60874 189922 60970 189978
rect 61026 189922 61094 189978
rect 61150 189922 61218 189978
rect 61274 189922 61342 189978
rect 61398 189922 61494 189978
rect 60874 172350 61494 189922
rect 69808 190350 70128 190384
rect 69808 190294 69878 190350
rect 69934 190294 70002 190350
rect 70058 190294 70128 190350
rect 69808 190226 70128 190294
rect 69808 190170 69878 190226
rect 69934 190170 70002 190226
rect 70058 190170 70128 190226
rect 69808 190102 70128 190170
rect 69808 190046 69878 190102
rect 69934 190046 70002 190102
rect 70058 190046 70128 190102
rect 69808 189978 70128 190046
rect 69808 189922 69878 189978
rect 69934 189922 70002 189978
rect 70058 189922 70128 189978
rect 69808 189888 70128 189922
rect 75154 184350 75774 201922
rect 75154 184294 75250 184350
rect 75306 184294 75374 184350
rect 75430 184294 75498 184350
rect 75554 184294 75622 184350
rect 75678 184294 75774 184350
rect 75154 184226 75774 184294
rect 75154 184170 75250 184226
rect 75306 184170 75374 184226
rect 75430 184170 75498 184226
rect 75554 184170 75622 184226
rect 75678 184170 75774 184226
rect 75154 184102 75774 184170
rect 75154 184046 75250 184102
rect 75306 184046 75374 184102
rect 75430 184046 75498 184102
rect 75554 184046 75622 184102
rect 75678 184046 75774 184102
rect 75154 183978 75774 184046
rect 75154 183922 75250 183978
rect 75306 183922 75374 183978
rect 75430 183922 75498 183978
rect 75554 183922 75622 183978
rect 75678 183922 75774 183978
rect 60874 172294 60970 172350
rect 61026 172294 61094 172350
rect 61150 172294 61218 172350
rect 61274 172294 61342 172350
rect 61398 172294 61494 172350
rect 60874 172226 61494 172294
rect 60874 172170 60970 172226
rect 61026 172170 61094 172226
rect 61150 172170 61218 172226
rect 61274 172170 61342 172226
rect 61398 172170 61494 172226
rect 60874 172102 61494 172170
rect 60874 172046 60970 172102
rect 61026 172046 61094 172102
rect 61150 172046 61218 172102
rect 61274 172046 61342 172102
rect 61398 172046 61494 172102
rect 60874 171978 61494 172046
rect 60874 171922 60970 171978
rect 61026 171922 61094 171978
rect 61150 171922 61218 171978
rect 61274 171922 61342 171978
rect 61398 171922 61494 171978
rect 60874 154350 61494 171922
rect 69808 172350 70128 172384
rect 69808 172294 69878 172350
rect 69934 172294 70002 172350
rect 70058 172294 70128 172350
rect 69808 172226 70128 172294
rect 69808 172170 69878 172226
rect 69934 172170 70002 172226
rect 70058 172170 70128 172226
rect 69808 172102 70128 172170
rect 69808 172046 69878 172102
rect 69934 172046 70002 172102
rect 70058 172046 70128 172102
rect 69808 171978 70128 172046
rect 69808 171922 69878 171978
rect 69934 171922 70002 171978
rect 70058 171922 70128 171978
rect 69808 171888 70128 171922
rect 75154 166350 75774 183922
rect 75154 166294 75250 166350
rect 75306 166294 75374 166350
rect 75430 166294 75498 166350
rect 75554 166294 75622 166350
rect 75678 166294 75774 166350
rect 75154 166226 75774 166294
rect 75154 166170 75250 166226
rect 75306 166170 75374 166226
rect 75430 166170 75498 166226
rect 75554 166170 75622 166226
rect 75678 166170 75774 166226
rect 75154 166102 75774 166170
rect 75154 166046 75250 166102
rect 75306 166046 75374 166102
rect 75430 166046 75498 166102
rect 75554 166046 75622 166102
rect 75678 166046 75774 166102
rect 75154 165978 75774 166046
rect 75154 165922 75250 165978
rect 75306 165922 75374 165978
rect 75430 165922 75498 165978
rect 75554 165922 75622 165978
rect 75678 165922 75774 165978
rect 60874 154294 60970 154350
rect 61026 154294 61094 154350
rect 61150 154294 61218 154350
rect 61274 154294 61342 154350
rect 61398 154294 61494 154350
rect 60874 154226 61494 154294
rect 60874 154170 60970 154226
rect 61026 154170 61094 154226
rect 61150 154170 61218 154226
rect 61274 154170 61342 154226
rect 61398 154170 61494 154226
rect 60874 154102 61494 154170
rect 60874 154046 60970 154102
rect 61026 154046 61094 154102
rect 61150 154046 61218 154102
rect 61274 154046 61342 154102
rect 61398 154046 61494 154102
rect 60874 153978 61494 154046
rect 60874 153922 60970 153978
rect 61026 153922 61094 153978
rect 61150 153922 61218 153978
rect 61274 153922 61342 153978
rect 61398 153922 61494 153978
rect 60874 136350 61494 153922
rect 69808 154350 70128 154384
rect 69808 154294 69878 154350
rect 69934 154294 70002 154350
rect 70058 154294 70128 154350
rect 69808 154226 70128 154294
rect 69808 154170 69878 154226
rect 69934 154170 70002 154226
rect 70058 154170 70128 154226
rect 69808 154102 70128 154170
rect 69808 154046 69878 154102
rect 69934 154046 70002 154102
rect 70058 154046 70128 154102
rect 69808 153978 70128 154046
rect 69808 153922 69878 153978
rect 69934 153922 70002 153978
rect 70058 153922 70128 153978
rect 69808 153888 70128 153922
rect 75154 148350 75774 165922
rect 75154 148294 75250 148350
rect 75306 148294 75374 148350
rect 75430 148294 75498 148350
rect 75554 148294 75622 148350
rect 75678 148294 75774 148350
rect 75154 148226 75774 148294
rect 75154 148170 75250 148226
rect 75306 148170 75374 148226
rect 75430 148170 75498 148226
rect 75554 148170 75622 148226
rect 75678 148170 75774 148226
rect 75154 148102 75774 148170
rect 75154 148046 75250 148102
rect 75306 148046 75374 148102
rect 75430 148046 75498 148102
rect 75554 148046 75622 148102
rect 75678 148046 75774 148102
rect 75154 147978 75774 148046
rect 75154 147922 75250 147978
rect 75306 147922 75374 147978
rect 75430 147922 75498 147978
rect 75554 147922 75622 147978
rect 75678 147922 75774 147978
rect 60874 136294 60970 136350
rect 61026 136294 61094 136350
rect 61150 136294 61218 136350
rect 61274 136294 61342 136350
rect 61398 136294 61494 136350
rect 60874 136226 61494 136294
rect 60874 136170 60970 136226
rect 61026 136170 61094 136226
rect 61150 136170 61218 136226
rect 61274 136170 61342 136226
rect 61398 136170 61494 136226
rect 60874 136102 61494 136170
rect 60874 136046 60970 136102
rect 61026 136046 61094 136102
rect 61150 136046 61218 136102
rect 61274 136046 61342 136102
rect 61398 136046 61494 136102
rect 60874 135978 61494 136046
rect 60874 135922 60970 135978
rect 61026 135922 61094 135978
rect 61150 135922 61218 135978
rect 61274 135922 61342 135978
rect 61398 135922 61494 135978
rect 60874 118350 61494 135922
rect 69808 136350 70128 136384
rect 69808 136294 69878 136350
rect 69934 136294 70002 136350
rect 70058 136294 70128 136350
rect 69808 136226 70128 136294
rect 69808 136170 69878 136226
rect 69934 136170 70002 136226
rect 70058 136170 70128 136226
rect 69808 136102 70128 136170
rect 69808 136046 69878 136102
rect 69934 136046 70002 136102
rect 70058 136046 70128 136102
rect 69808 135978 70128 136046
rect 69808 135922 69878 135978
rect 69934 135922 70002 135978
rect 70058 135922 70128 135978
rect 69808 135888 70128 135922
rect 75154 130350 75774 147922
rect 75154 130294 75250 130350
rect 75306 130294 75374 130350
rect 75430 130294 75498 130350
rect 75554 130294 75622 130350
rect 75678 130294 75774 130350
rect 75154 130226 75774 130294
rect 75154 130170 75250 130226
rect 75306 130170 75374 130226
rect 75430 130170 75498 130226
rect 75554 130170 75622 130226
rect 75678 130170 75774 130226
rect 75154 130102 75774 130170
rect 75154 130046 75250 130102
rect 75306 130046 75374 130102
rect 75430 130046 75498 130102
rect 75554 130046 75622 130102
rect 75678 130046 75774 130102
rect 75154 129978 75774 130046
rect 75154 129922 75250 129978
rect 75306 129922 75374 129978
rect 75430 129922 75498 129978
rect 75554 129922 75622 129978
rect 75678 129922 75774 129978
rect 60874 118294 60970 118350
rect 61026 118294 61094 118350
rect 61150 118294 61218 118350
rect 61274 118294 61342 118350
rect 61398 118294 61494 118350
rect 60874 118226 61494 118294
rect 60874 118170 60970 118226
rect 61026 118170 61094 118226
rect 61150 118170 61218 118226
rect 61274 118170 61342 118226
rect 61398 118170 61494 118226
rect 60874 118102 61494 118170
rect 60874 118046 60970 118102
rect 61026 118046 61094 118102
rect 61150 118046 61218 118102
rect 61274 118046 61342 118102
rect 61398 118046 61494 118102
rect 60874 117978 61494 118046
rect 60874 117922 60970 117978
rect 61026 117922 61094 117978
rect 61150 117922 61218 117978
rect 61274 117922 61342 117978
rect 61398 117922 61494 117978
rect 60874 100350 61494 117922
rect 69808 118350 70128 118384
rect 69808 118294 69878 118350
rect 69934 118294 70002 118350
rect 70058 118294 70128 118350
rect 69808 118226 70128 118294
rect 69808 118170 69878 118226
rect 69934 118170 70002 118226
rect 70058 118170 70128 118226
rect 69808 118102 70128 118170
rect 69808 118046 69878 118102
rect 69934 118046 70002 118102
rect 70058 118046 70128 118102
rect 69808 117978 70128 118046
rect 69808 117922 69878 117978
rect 69934 117922 70002 117978
rect 70058 117922 70128 117978
rect 69808 117888 70128 117922
rect 75154 112350 75774 129922
rect 75154 112294 75250 112350
rect 75306 112294 75374 112350
rect 75430 112294 75498 112350
rect 75554 112294 75622 112350
rect 75678 112294 75774 112350
rect 75154 112226 75774 112294
rect 75154 112170 75250 112226
rect 75306 112170 75374 112226
rect 75430 112170 75498 112226
rect 75554 112170 75622 112226
rect 75678 112170 75774 112226
rect 75154 112102 75774 112170
rect 75154 112046 75250 112102
rect 75306 112046 75374 112102
rect 75430 112046 75498 112102
rect 75554 112046 75622 112102
rect 75678 112046 75774 112102
rect 75154 111978 75774 112046
rect 75154 111922 75250 111978
rect 75306 111922 75374 111978
rect 75430 111922 75498 111978
rect 75554 111922 75622 111978
rect 75678 111922 75774 111978
rect 60874 100294 60970 100350
rect 61026 100294 61094 100350
rect 61150 100294 61218 100350
rect 61274 100294 61342 100350
rect 61398 100294 61494 100350
rect 60874 100226 61494 100294
rect 60874 100170 60970 100226
rect 61026 100170 61094 100226
rect 61150 100170 61218 100226
rect 61274 100170 61342 100226
rect 61398 100170 61494 100226
rect 60874 100102 61494 100170
rect 60874 100046 60970 100102
rect 61026 100046 61094 100102
rect 61150 100046 61218 100102
rect 61274 100046 61342 100102
rect 61398 100046 61494 100102
rect 60874 99978 61494 100046
rect 60874 99922 60970 99978
rect 61026 99922 61094 99978
rect 61150 99922 61218 99978
rect 61274 99922 61342 99978
rect 61398 99922 61494 99978
rect 60874 82350 61494 99922
rect 69808 100350 70128 100384
rect 69808 100294 69878 100350
rect 69934 100294 70002 100350
rect 70058 100294 70128 100350
rect 69808 100226 70128 100294
rect 69808 100170 69878 100226
rect 69934 100170 70002 100226
rect 70058 100170 70128 100226
rect 69808 100102 70128 100170
rect 69808 100046 69878 100102
rect 69934 100046 70002 100102
rect 70058 100046 70128 100102
rect 69808 99978 70128 100046
rect 69808 99922 69878 99978
rect 69934 99922 70002 99978
rect 70058 99922 70128 99978
rect 69808 99888 70128 99922
rect 75154 94350 75774 111922
rect 75154 94294 75250 94350
rect 75306 94294 75374 94350
rect 75430 94294 75498 94350
rect 75554 94294 75622 94350
rect 75678 94294 75774 94350
rect 75154 94226 75774 94294
rect 75154 94170 75250 94226
rect 75306 94170 75374 94226
rect 75430 94170 75498 94226
rect 75554 94170 75622 94226
rect 75678 94170 75774 94226
rect 75154 94102 75774 94170
rect 75154 94046 75250 94102
rect 75306 94046 75374 94102
rect 75430 94046 75498 94102
rect 75554 94046 75622 94102
rect 75678 94046 75774 94102
rect 75154 93978 75774 94046
rect 75154 93922 75250 93978
rect 75306 93922 75374 93978
rect 75430 93922 75498 93978
rect 75554 93922 75622 93978
rect 75678 93922 75774 93978
rect 60874 82294 60970 82350
rect 61026 82294 61094 82350
rect 61150 82294 61218 82350
rect 61274 82294 61342 82350
rect 61398 82294 61494 82350
rect 60874 82226 61494 82294
rect 60874 82170 60970 82226
rect 61026 82170 61094 82226
rect 61150 82170 61218 82226
rect 61274 82170 61342 82226
rect 61398 82170 61494 82226
rect 60874 82102 61494 82170
rect 60874 82046 60970 82102
rect 61026 82046 61094 82102
rect 61150 82046 61218 82102
rect 61274 82046 61342 82102
rect 61398 82046 61494 82102
rect 60874 81978 61494 82046
rect 60874 81922 60970 81978
rect 61026 81922 61094 81978
rect 61150 81922 61218 81978
rect 61274 81922 61342 81978
rect 61398 81922 61494 81978
rect 60874 64350 61494 81922
rect 69808 82350 70128 82384
rect 69808 82294 69878 82350
rect 69934 82294 70002 82350
rect 70058 82294 70128 82350
rect 69808 82226 70128 82294
rect 69808 82170 69878 82226
rect 69934 82170 70002 82226
rect 70058 82170 70128 82226
rect 69808 82102 70128 82170
rect 69808 82046 69878 82102
rect 69934 82046 70002 82102
rect 70058 82046 70128 82102
rect 69808 81978 70128 82046
rect 69808 81922 69878 81978
rect 69934 81922 70002 81978
rect 70058 81922 70128 81978
rect 69808 81888 70128 81922
rect 75154 76350 75774 93922
rect 75154 76294 75250 76350
rect 75306 76294 75374 76350
rect 75430 76294 75498 76350
rect 75554 76294 75622 76350
rect 75678 76294 75774 76350
rect 75154 76226 75774 76294
rect 75154 76170 75250 76226
rect 75306 76170 75374 76226
rect 75430 76170 75498 76226
rect 75554 76170 75622 76226
rect 75678 76170 75774 76226
rect 75154 76102 75774 76170
rect 75154 76046 75250 76102
rect 75306 76046 75374 76102
rect 75430 76046 75498 76102
rect 75554 76046 75622 76102
rect 75678 76046 75774 76102
rect 75154 75978 75774 76046
rect 75154 75922 75250 75978
rect 75306 75922 75374 75978
rect 75430 75922 75498 75978
rect 75554 75922 75622 75978
rect 75678 75922 75774 75978
rect 60874 64294 60970 64350
rect 61026 64294 61094 64350
rect 61150 64294 61218 64350
rect 61274 64294 61342 64350
rect 61398 64294 61494 64350
rect 60874 64226 61494 64294
rect 60874 64170 60970 64226
rect 61026 64170 61094 64226
rect 61150 64170 61218 64226
rect 61274 64170 61342 64226
rect 61398 64170 61494 64226
rect 60874 64102 61494 64170
rect 60874 64046 60970 64102
rect 61026 64046 61094 64102
rect 61150 64046 61218 64102
rect 61274 64046 61342 64102
rect 61398 64046 61494 64102
rect 60874 63978 61494 64046
rect 60874 63922 60970 63978
rect 61026 63922 61094 63978
rect 61150 63922 61218 63978
rect 61274 63922 61342 63978
rect 61398 63922 61494 63978
rect 60874 46350 61494 63922
rect 69808 64350 70128 64384
rect 69808 64294 69878 64350
rect 69934 64294 70002 64350
rect 70058 64294 70128 64350
rect 69808 64226 70128 64294
rect 69808 64170 69878 64226
rect 69934 64170 70002 64226
rect 70058 64170 70128 64226
rect 69808 64102 70128 64170
rect 69808 64046 69878 64102
rect 69934 64046 70002 64102
rect 70058 64046 70128 64102
rect 69808 63978 70128 64046
rect 69808 63922 69878 63978
rect 69934 63922 70002 63978
rect 70058 63922 70128 63978
rect 69808 63888 70128 63922
rect 75154 58350 75774 75922
rect 75154 58294 75250 58350
rect 75306 58294 75374 58350
rect 75430 58294 75498 58350
rect 75554 58294 75622 58350
rect 75678 58294 75774 58350
rect 75154 58226 75774 58294
rect 75154 58170 75250 58226
rect 75306 58170 75374 58226
rect 75430 58170 75498 58226
rect 75554 58170 75622 58226
rect 75678 58170 75774 58226
rect 75154 58102 75774 58170
rect 75154 58046 75250 58102
rect 75306 58046 75374 58102
rect 75430 58046 75498 58102
rect 75554 58046 75622 58102
rect 75678 58046 75774 58102
rect 75154 57978 75774 58046
rect 75154 57922 75250 57978
rect 75306 57922 75374 57978
rect 75430 57922 75498 57978
rect 75554 57922 75622 57978
rect 75678 57922 75774 57978
rect 60874 46294 60970 46350
rect 61026 46294 61094 46350
rect 61150 46294 61218 46350
rect 61274 46294 61342 46350
rect 61398 46294 61494 46350
rect 60874 46226 61494 46294
rect 60874 46170 60970 46226
rect 61026 46170 61094 46226
rect 61150 46170 61218 46226
rect 61274 46170 61342 46226
rect 61398 46170 61494 46226
rect 60874 46102 61494 46170
rect 60874 46046 60970 46102
rect 61026 46046 61094 46102
rect 61150 46046 61218 46102
rect 61274 46046 61342 46102
rect 61398 46046 61494 46102
rect 60874 45978 61494 46046
rect 60874 45922 60970 45978
rect 61026 45922 61094 45978
rect 61150 45922 61218 45978
rect 61274 45922 61342 45978
rect 61398 45922 61494 45978
rect 60874 28350 61494 45922
rect 69808 46350 70128 46384
rect 69808 46294 69878 46350
rect 69934 46294 70002 46350
rect 70058 46294 70128 46350
rect 69808 46226 70128 46294
rect 69808 46170 69878 46226
rect 69934 46170 70002 46226
rect 70058 46170 70128 46226
rect 69808 46102 70128 46170
rect 69808 46046 69878 46102
rect 69934 46046 70002 46102
rect 70058 46046 70128 46102
rect 69808 45978 70128 46046
rect 69808 45922 69878 45978
rect 69934 45922 70002 45978
rect 70058 45922 70128 45978
rect 69808 45888 70128 45922
rect 60874 28294 60970 28350
rect 61026 28294 61094 28350
rect 61150 28294 61218 28350
rect 61274 28294 61342 28350
rect 61398 28294 61494 28350
rect 60874 28226 61494 28294
rect 60874 28170 60970 28226
rect 61026 28170 61094 28226
rect 61150 28170 61218 28226
rect 61274 28170 61342 28226
rect 61398 28170 61494 28226
rect 60874 28102 61494 28170
rect 60874 28046 60970 28102
rect 61026 28046 61094 28102
rect 61150 28046 61218 28102
rect 61274 28046 61342 28102
rect 61398 28046 61494 28102
rect 60874 27978 61494 28046
rect 60874 27922 60970 27978
rect 61026 27922 61094 27978
rect 61150 27922 61218 27978
rect 61274 27922 61342 27978
rect 61398 27922 61494 27978
rect 60874 10350 61494 27922
rect 60874 10294 60970 10350
rect 61026 10294 61094 10350
rect 61150 10294 61218 10350
rect 61274 10294 61342 10350
rect 61398 10294 61494 10350
rect 60874 10226 61494 10294
rect 60874 10170 60970 10226
rect 61026 10170 61094 10226
rect 61150 10170 61218 10226
rect 61274 10170 61342 10226
rect 61398 10170 61494 10226
rect 60874 10102 61494 10170
rect 60874 10046 60970 10102
rect 61026 10046 61094 10102
rect 61150 10046 61218 10102
rect 61274 10046 61342 10102
rect 61398 10046 61494 10102
rect 60874 9978 61494 10046
rect 60874 9922 60970 9978
rect 61026 9922 61094 9978
rect 61150 9922 61218 9978
rect 61274 9922 61342 9978
rect 61398 9922 61494 9978
rect 60874 -1120 61494 9922
rect 60874 -1176 60970 -1120
rect 61026 -1176 61094 -1120
rect 61150 -1176 61218 -1120
rect 61274 -1176 61342 -1120
rect 61398 -1176 61494 -1120
rect 60874 -1244 61494 -1176
rect 60874 -1300 60970 -1244
rect 61026 -1300 61094 -1244
rect 61150 -1300 61218 -1244
rect 61274 -1300 61342 -1244
rect 61398 -1300 61494 -1244
rect 60874 -1368 61494 -1300
rect 60874 -1424 60970 -1368
rect 61026 -1424 61094 -1368
rect 61150 -1424 61218 -1368
rect 61274 -1424 61342 -1368
rect 61398 -1424 61494 -1368
rect 60874 -1492 61494 -1424
rect 60874 -1548 60970 -1492
rect 61026 -1548 61094 -1492
rect 61150 -1548 61218 -1492
rect 61274 -1548 61342 -1492
rect 61398 -1548 61494 -1492
rect 60874 -1644 61494 -1548
rect 75154 40350 75774 57922
rect 75154 40294 75250 40350
rect 75306 40294 75374 40350
rect 75430 40294 75498 40350
rect 75554 40294 75622 40350
rect 75678 40294 75774 40350
rect 75154 40226 75774 40294
rect 75154 40170 75250 40226
rect 75306 40170 75374 40226
rect 75430 40170 75498 40226
rect 75554 40170 75622 40226
rect 75678 40170 75774 40226
rect 75154 40102 75774 40170
rect 75154 40046 75250 40102
rect 75306 40046 75374 40102
rect 75430 40046 75498 40102
rect 75554 40046 75622 40102
rect 75678 40046 75774 40102
rect 75154 39978 75774 40046
rect 75154 39922 75250 39978
rect 75306 39922 75374 39978
rect 75430 39922 75498 39978
rect 75554 39922 75622 39978
rect 75678 39922 75774 39978
rect 75154 22350 75774 39922
rect 75154 22294 75250 22350
rect 75306 22294 75374 22350
rect 75430 22294 75498 22350
rect 75554 22294 75622 22350
rect 75678 22294 75774 22350
rect 75154 22226 75774 22294
rect 75154 22170 75250 22226
rect 75306 22170 75374 22226
rect 75430 22170 75498 22226
rect 75554 22170 75622 22226
rect 75678 22170 75774 22226
rect 75154 22102 75774 22170
rect 75154 22046 75250 22102
rect 75306 22046 75374 22102
rect 75430 22046 75498 22102
rect 75554 22046 75622 22102
rect 75678 22046 75774 22102
rect 75154 21978 75774 22046
rect 75154 21922 75250 21978
rect 75306 21922 75374 21978
rect 75430 21922 75498 21978
rect 75554 21922 75622 21978
rect 75678 21922 75774 21978
rect 75154 4350 75774 21922
rect 75154 4294 75250 4350
rect 75306 4294 75374 4350
rect 75430 4294 75498 4350
rect 75554 4294 75622 4350
rect 75678 4294 75774 4350
rect 75154 4226 75774 4294
rect 75154 4170 75250 4226
rect 75306 4170 75374 4226
rect 75430 4170 75498 4226
rect 75554 4170 75622 4226
rect 75678 4170 75774 4226
rect 75154 4102 75774 4170
rect 75154 4046 75250 4102
rect 75306 4046 75374 4102
rect 75430 4046 75498 4102
rect 75554 4046 75622 4102
rect 75678 4046 75774 4102
rect 75154 3978 75774 4046
rect 75154 3922 75250 3978
rect 75306 3922 75374 3978
rect 75430 3922 75498 3978
rect 75554 3922 75622 3978
rect 75678 3922 75774 3978
rect 75154 -160 75774 3922
rect 75154 -216 75250 -160
rect 75306 -216 75374 -160
rect 75430 -216 75498 -160
rect 75554 -216 75622 -160
rect 75678 -216 75774 -160
rect 75154 -284 75774 -216
rect 75154 -340 75250 -284
rect 75306 -340 75374 -284
rect 75430 -340 75498 -284
rect 75554 -340 75622 -284
rect 75678 -340 75774 -284
rect 75154 -408 75774 -340
rect 75154 -464 75250 -408
rect 75306 -464 75374 -408
rect 75430 -464 75498 -408
rect 75554 -464 75622 -408
rect 75678 -464 75774 -408
rect 75154 -532 75774 -464
rect 75154 -588 75250 -532
rect 75306 -588 75374 -532
rect 75430 -588 75498 -532
rect 75554 -588 75622 -532
rect 75678 -588 75774 -532
rect 75154 -1644 75774 -588
rect 78874 598172 79494 598268
rect 78874 598116 78970 598172
rect 79026 598116 79094 598172
rect 79150 598116 79218 598172
rect 79274 598116 79342 598172
rect 79398 598116 79494 598172
rect 78874 598048 79494 598116
rect 78874 597992 78970 598048
rect 79026 597992 79094 598048
rect 79150 597992 79218 598048
rect 79274 597992 79342 598048
rect 79398 597992 79494 598048
rect 78874 597924 79494 597992
rect 78874 597868 78970 597924
rect 79026 597868 79094 597924
rect 79150 597868 79218 597924
rect 79274 597868 79342 597924
rect 79398 597868 79494 597924
rect 78874 597800 79494 597868
rect 78874 597744 78970 597800
rect 79026 597744 79094 597800
rect 79150 597744 79218 597800
rect 79274 597744 79342 597800
rect 79398 597744 79494 597800
rect 78874 586350 79494 597744
rect 78874 586294 78970 586350
rect 79026 586294 79094 586350
rect 79150 586294 79218 586350
rect 79274 586294 79342 586350
rect 79398 586294 79494 586350
rect 78874 586226 79494 586294
rect 78874 586170 78970 586226
rect 79026 586170 79094 586226
rect 79150 586170 79218 586226
rect 79274 586170 79342 586226
rect 79398 586170 79494 586226
rect 78874 586102 79494 586170
rect 78874 586046 78970 586102
rect 79026 586046 79094 586102
rect 79150 586046 79218 586102
rect 79274 586046 79342 586102
rect 79398 586046 79494 586102
rect 78874 585978 79494 586046
rect 78874 585922 78970 585978
rect 79026 585922 79094 585978
rect 79150 585922 79218 585978
rect 79274 585922 79342 585978
rect 79398 585922 79494 585978
rect 78874 568350 79494 585922
rect 78874 568294 78970 568350
rect 79026 568294 79094 568350
rect 79150 568294 79218 568350
rect 79274 568294 79342 568350
rect 79398 568294 79494 568350
rect 78874 568226 79494 568294
rect 78874 568170 78970 568226
rect 79026 568170 79094 568226
rect 79150 568170 79218 568226
rect 79274 568170 79342 568226
rect 79398 568170 79494 568226
rect 78874 568102 79494 568170
rect 78874 568046 78970 568102
rect 79026 568046 79094 568102
rect 79150 568046 79218 568102
rect 79274 568046 79342 568102
rect 79398 568046 79494 568102
rect 78874 567978 79494 568046
rect 78874 567922 78970 567978
rect 79026 567922 79094 567978
rect 79150 567922 79218 567978
rect 79274 567922 79342 567978
rect 79398 567922 79494 567978
rect 78874 550350 79494 567922
rect 78874 550294 78970 550350
rect 79026 550294 79094 550350
rect 79150 550294 79218 550350
rect 79274 550294 79342 550350
rect 79398 550294 79494 550350
rect 78874 550226 79494 550294
rect 78874 550170 78970 550226
rect 79026 550170 79094 550226
rect 79150 550170 79218 550226
rect 79274 550170 79342 550226
rect 79398 550170 79494 550226
rect 78874 550102 79494 550170
rect 78874 550046 78970 550102
rect 79026 550046 79094 550102
rect 79150 550046 79218 550102
rect 79274 550046 79342 550102
rect 79398 550046 79494 550102
rect 78874 549978 79494 550046
rect 78874 549922 78970 549978
rect 79026 549922 79094 549978
rect 79150 549922 79218 549978
rect 79274 549922 79342 549978
rect 79398 549922 79494 549978
rect 78874 532350 79494 549922
rect 78874 532294 78970 532350
rect 79026 532294 79094 532350
rect 79150 532294 79218 532350
rect 79274 532294 79342 532350
rect 79398 532294 79494 532350
rect 78874 532226 79494 532294
rect 78874 532170 78970 532226
rect 79026 532170 79094 532226
rect 79150 532170 79218 532226
rect 79274 532170 79342 532226
rect 79398 532170 79494 532226
rect 78874 532102 79494 532170
rect 78874 532046 78970 532102
rect 79026 532046 79094 532102
rect 79150 532046 79218 532102
rect 79274 532046 79342 532102
rect 79398 532046 79494 532102
rect 78874 531978 79494 532046
rect 78874 531922 78970 531978
rect 79026 531922 79094 531978
rect 79150 531922 79218 531978
rect 79274 531922 79342 531978
rect 79398 531922 79494 531978
rect 78874 514350 79494 531922
rect 93154 597212 93774 598268
rect 93154 597156 93250 597212
rect 93306 597156 93374 597212
rect 93430 597156 93498 597212
rect 93554 597156 93622 597212
rect 93678 597156 93774 597212
rect 93154 597088 93774 597156
rect 93154 597032 93250 597088
rect 93306 597032 93374 597088
rect 93430 597032 93498 597088
rect 93554 597032 93622 597088
rect 93678 597032 93774 597088
rect 93154 596964 93774 597032
rect 93154 596908 93250 596964
rect 93306 596908 93374 596964
rect 93430 596908 93498 596964
rect 93554 596908 93622 596964
rect 93678 596908 93774 596964
rect 93154 596840 93774 596908
rect 93154 596784 93250 596840
rect 93306 596784 93374 596840
rect 93430 596784 93498 596840
rect 93554 596784 93622 596840
rect 93678 596784 93774 596840
rect 93154 580350 93774 596784
rect 93154 580294 93250 580350
rect 93306 580294 93374 580350
rect 93430 580294 93498 580350
rect 93554 580294 93622 580350
rect 93678 580294 93774 580350
rect 93154 580226 93774 580294
rect 93154 580170 93250 580226
rect 93306 580170 93374 580226
rect 93430 580170 93498 580226
rect 93554 580170 93622 580226
rect 93678 580170 93774 580226
rect 93154 580102 93774 580170
rect 93154 580046 93250 580102
rect 93306 580046 93374 580102
rect 93430 580046 93498 580102
rect 93554 580046 93622 580102
rect 93678 580046 93774 580102
rect 93154 579978 93774 580046
rect 93154 579922 93250 579978
rect 93306 579922 93374 579978
rect 93430 579922 93498 579978
rect 93554 579922 93622 579978
rect 93678 579922 93774 579978
rect 93154 562350 93774 579922
rect 93154 562294 93250 562350
rect 93306 562294 93374 562350
rect 93430 562294 93498 562350
rect 93554 562294 93622 562350
rect 93678 562294 93774 562350
rect 93154 562226 93774 562294
rect 93154 562170 93250 562226
rect 93306 562170 93374 562226
rect 93430 562170 93498 562226
rect 93554 562170 93622 562226
rect 93678 562170 93774 562226
rect 93154 562102 93774 562170
rect 93154 562046 93250 562102
rect 93306 562046 93374 562102
rect 93430 562046 93498 562102
rect 93554 562046 93622 562102
rect 93678 562046 93774 562102
rect 93154 561978 93774 562046
rect 93154 561922 93250 561978
rect 93306 561922 93374 561978
rect 93430 561922 93498 561978
rect 93554 561922 93622 561978
rect 93678 561922 93774 561978
rect 93154 544350 93774 561922
rect 93154 544294 93250 544350
rect 93306 544294 93374 544350
rect 93430 544294 93498 544350
rect 93554 544294 93622 544350
rect 93678 544294 93774 544350
rect 93154 544226 93774 544294
rect 93154 544170 93250 544226
rect 93306 544170 93374 544226
rect 93430 544170 93498 544226
rect 93554 544170 93622 544226
rect 93678 544170 93774 544226
rect 93154 544102 93774 544170
rect 93154 544046 93250 544102
rect 93306 544046 93374 544102
rect 93430 544046 93498 544102
rect 93554 544046 93622 544102
rect 93678 544046 93774 544102
rect 93154 543978 93774 544046
rect 93154 543922 93250 543978
rect 93306 543922 93374 543978
rect 93430 543922 93498 543978
rect 93554 543922 93622 543978
rect 93678 543922 93774 543978
rect 93154 526350 93774 543922
rect 85168 526293 85488 526332
rect 85168 526237 85238 526293
rect 85294 526237 85362 526293
rect 85418 526237 85488 526293
rect 85168 526169 85488 526237
rect 85168 526113 85238 526169
rect 85294 526113 85362 526169
rect 85418 526113 85488 526169
rect 85168 526045 85488 526113
rect 85168 525989 85238 526045
rect 85294 525989 85362 526045
rect 85418 525989 85488 526045
rect 85168 525921 85488 525989
rect 85168 525865 85238 525921
rect 85294 525865 85362 525921
rect 85418 525865 85488 525921
rect 85168 525826 85488 525865
rect 93154 526294 93250 526350
rect 93306 526294 93374 526350
rect 93430 526294 93498 526350
rect 93554 526294 93622 526350
rect 93678 526294 93774 526350
rect 93154 526226 93774 526294
rect 93154 526170 93250 526226
rect 93306 526170 93374 526226
rect 93430 526170 93498 526226
rect 93554 526170 93622 526226
rect 93678 526170 93774 526226
rect 93154 526102 93774 526170
rect 93154 526046 93250 526102
rect 93306 526046 93374 526102
rect 93430 526046 93498 526102
rect 93554 526046 93622 526102
rect 93678 526046 93774 526102
rect 93154 525978 93774 526046
rect 93154 525922 93250 525978
rect 93306 525922 93374 525978
rect 93430 525922 93498 525978
rect 93554 525922 93622 525978
rect 93678 525922 93774 525978
rect 78874 514294 78970 514350
rect 79026 514294 79094 514350
rect 79150 514294 79218 514350
rect 79274 514294 79342 514350
rect 79398 514294 79494 514350
rect 78874 514226 79494 514294
rect 78874 514170 78970 514226
rect 79026 514170 79094 514226
rect 79150 514170 79218 514226
rect 79274 514170 79342 514226
rect 79398 514170 79494 514226
rect 78874 514102 79494 514170
rect 78874 514046 78970 514102
rect 79026 514046 79094 514102
rect 79150 514046 79218 514102
rect 79274 514046 79342 514102
rect 79398 514046 79494 514102
rect 78874 513978 79494 514046
rect 78874 513922 78970 513978
rect 79026 513922 79094 513978
rect 79150 513922 79218 513978
rect 79274 513922 79342 513978
rect 79398 513922 79494 513978
rect 78874 496350 79494 513922
rect 85168 508350 85488 508384
rect 85168 508294 85238 508350
rect 85294 508294 85362 508350
rect 85418 508294 85488 508350
rect 85168 508226 85488 508294
rect 85168 508170 85238 508226
rect 85294 508170 85362 508226
rect 85418 508170 85488 508226
rect 85168 508102 85488 508170
rect 85168 508046 85238 508102
rect 85294 508046 85362 508102
rect 85418 508046 85488 508102
rect 85168 507978 85488 508046
rect 85168 507922 85238 507978
rect 85294 507922 85362 507978
rect 85418 507922 85488 507978
rect 85168 507888 85488 507922
rect 93154 508350 93774 525922
rect 93154 508294 93250 508350
rect 93306 508294 93374 508350
rect 93430 508294 93498 508350
rect 93554 508294 93622 508350
rect 93678 508294 93774 508350
rect 93154 508226 93774 508294
rect 93154 508170 93250 508226
rect 93306 508170 93374 508226
rect 93430 508170 93498 508226
rect 93554 508170 93622 508226
rect 93678 508170 93774 508226
rect 93154 508102 93774 508170
rect 93154 508046 93250 508102
rect 93306 508046 93374 508102
rect 93430 508046 93498 508102
rect 93554 508046 93622 508102
rect 93678 508046 93774 508102
rect 93154 507978 93774 508046
rect 93154 507922 93250 507978
rect 93306 507922 93374 507978
rect 93430 507922 93498 507978
rect 93554 507922 93622 507978
rect 93678 507922 93774 507978
rect 78874 496294 78970 496350
rect 79026 496294 79094 496350
rect 79150 496294 79218 496350
rect 79274 496294 79342 496350
rect 79398 496294 79494 496350
rect 78874 496226 79494 496294
rect 78874 496170 78970 496226
rect 79026 496170 79094 496226
rect 79150 496170 79218 496226
rect 79274 496170 79342 496226
rect 79398 496170 79494 496226
rect 78874 496102 79494 496170
rect 78874 496046 78970 496102
rect 79026 496046 79094 496102
rect 79150 496046 79218 496102
rect 79274 496046 79342 496102
rect 79398 496046 79494 496102
rect 78874 495978 79494 496046
rect 78874 495922 78970 495978
rect 79026 495922 79094 495978
rect 79150 495922 79218 495978
rect 79274 495922 79342 495978
rect 79398 495922 79494 495978
rect 78874 478350 79494 495922
rect 85168 490350 85488 490384
rect 85168 490294 85238 490350
rect 85294 490294 85362 490350
rect 85418 490294 85488 490350
rect 85168 490226 85488 490294
rect 85168 490170 85238 490226
rect 85294 490170 85362 490226
rect 85418 490170 85488 490226
rect 85168 490102 85488 490170
rect 85168 490046 85238 490102
rect 85294 490046 85362 490102
rect 85418 490046 85488 490102
rect 85168 489978 85488 490046
rect 85168 489922 85238 489978
rect 85294 489922 85362 489978
rect 85418 489922 85488 489978
rect 85168 489888 85488 489922
rect 93154 490350 93774 507922
rect 93154 490294 93250 490350
rect 93306 490294 93374 490350
rect 93430 490294 93498 490350
rect 93554 490294 93622 490350
rect 93678 490294 93774 490350
rect 93154 490226 93774 490294
rect 93154 490170 93250 490226
rect 93306 490170 93374 490226
rect 93430 490170 93498 490226
rect 93554 490170 93622 490226
rect 93678 490170 93774 490226
rect 93154 490102 93774 490170
rect 93154 490046 93250 490102
rect 93306 490046 93374 490102
rect 93430 490046 93498 490102
rect 93554 490046 93622 490102
rect 93678 490046 93774 490102
rect 93154 489978 93774 490046
rect 93154 489922 93250 489978
rect 93306 489922 93374 489978
rect 93430 489922 93498 489978
rect 93554 489922 93622 489978
rect 93678 489922 93774 489978
rect 78874 478294 78970 478350
rect 79026 478294 79094 478350
rect 79150 478294 79218 478350
rect 79274 478294 79342 478350
rect 79398 478294 79494 478350
rect 78874 478226 79494 478294
rect 78874 478170 78970 478226
rect 79026 478170 79094 478226
rect 79150 478170 79218 478226
rect 79274 478170 79342 478226
rect 79398 478170 79494 478226
rect 78874 478102 79494 478170
rect 78874 478046 78970 478102
rect 79026 478046 79094 478102
rect 79150 478046 79218 478102
rect 79274 478046 79342 478102
rect 79398 478046 79494 478102
rect 78874 477978 79494 478046
rect 78874 477922 78970 477978
rect 79026 477922 79094 477978
rect 79150 477922 79218 477978
rect 79274 477922 79342 477978
rect 79398 477922 79494 477978
rect 78874 460350 79494 477922
rect 85168 472350 85488 472384
rect 85168 472294 85238 472350
rect 85294 472294 85362 472350
rect 85418 472294 85488 472350
rect 85168 472226 85488 472294
rect 85168 472170 85238 472226
rect 85294 472170 85362 472226
rect 85418 472170 85488 472226
rect 85168 472102 85488 472170
rect 85168 472046 85238 472102
rect 85294 472046 85362 472102
rect 85418 472046 85488 472102
rect 85168 471978 85488 472046
rect 85168 471922 85238 471978
rect 85294 471922 85362 471978
rect 85418 471922 85488 471978
rect 85168 471888 85488 471922
rect 93154 472350 93774 489922
rect 93154 472294 93250 472350
rect 93306 472294 93374 472350
rect 93430 472294 93498 472350
rect 93554 472294 93622 472350
rect 93678 472294 93774 472350
rect 93154 472226 93774 472294
rect 93154 472170 93250 472226
rect 93306 472170 93374 472226
rect 93430 472170 93498 472226
rect 93554 472170 93622 472226
rect 93678 472170 93774 472226
rect 93154 472102 93774 472170
rect 93154 472046 93250 472102
rect 93306 472046 93374 472102
rect 93430 472046 93498 472102
rect 93554 472046 93622 472102
rect 93678 472046 93774 472102
rect 93154 471978 93774 472046
rect 93154 471922 93250 471978
rect 93306 471922 93374 471978
rect 93430 471922 93498 471978
rect 93554 471922 93622 471978
rect 93678 471922 93774 471978
rect 78874 460294 78970 460350
rect 79026 460294 79094 460350
rect 79150 460294 79218 460350
rect 79274 460294 79342 460350
rect 79398 460294 79494 460350
rect 78874 460226 79494 460294
rect 78874 460170 78970 460226
rect 79026 460170 79094 460226
rect 79150 460170 79218 460226
rect 79274 460170 79342 460226
rect 79398 460170 79494 460226
rect 78874 460102 79494 460170
rect 78874 460046 78970 460102
rect 79026 460046 79094 460102
rect 79150 460046 79218 460102
rect 79274 460046 79342 460102
rect 79398 460046 79494 460102
rect 78874 459978 79494 460046
rect 78874 459922 78970 459978
rect 79026 459922 79094 459978
rect 79150 459922 79218 459978
rect 79274 459922 79342 459978
rect 79398 459922 79494 459978
rect 78874 442350 79494 459922
rect 85168 454350 85488 454384
rect 85168 454294 85238 454350
rect 85294 454294 85362 454350
rect 85418 454294 85488 454350
rect 85168 454226 85488 454294
rect 85168 454170 85238 454226
rect 85294 454170 85362 454226
rect 85418 454170 85488 454226
rect 85168 454102 85488 454170
rect 85168 454046 85238 454102
rect 85294 454046 85362 454102
rect 85418 454046 85488 454102
rect 85168 453978 85488 454046
rect 85168 453922 85238 453978
rect 85294 453922 85362 453978
rect 85418 453922 85488 453978
rect 85168 453888 85488 453922
rect 93154 454350 93774 471922
rect 93154 454294 93250 454350
rect 93306 454294 93374 454350
rect 93430 454294 93498 454350
rect 93554 454294 93622 454350
rect 93678 454294 93774 454350
rect 93154 454226 93774 454294
rect 93154 454170 93250 454226
rect 93306 454170 93374 454226
rect 93430 454170 93498 454226
rect 93554 454170 93622 454226
rect 93678 454170 93774 454226
rect 93154 454102 93774 454170
rect 93154 454046 93250 454102
rect 93306 454046 93374 454102
rect 93430 454046 93498 454102
rect 93554 454046 93622 454102
rect 93678 454046 93774 454102
rect 93154 453978 93774 454046
rect 93154 453922 93250 453978
rect 93306 453922 93374 453978
rect 93430 453922 93498 453978
rect 93554 453922 93622 453978
rect 93678 453922 93774 453978
rect 78874 442294 78970 442350
rect 79026 442294 79094 442350
rect 79150 442294 79218 442350
rect 79274 442294 79342 442350
rect 79398 442294 79494 442350
rect 78874 442226 79494 442294
rect 78874 442170 78970 442226
rect 79026 442170 79094 442226
rect 79150 442170 79218 442226
rect 79274 442170 79342 442226
rect 79398 442170 79494 442226
rect 78874 442102 79494 442170
rect 78874 442046 78970 442102
rect 79026 442046 79094 442102
rect 79150 442046 79218 442102
rect 79274 442046 79342 442102
rect 79398 442046 79494 442102
rect 78874 441978 79494 442046
rect 78874 441922 78970 441978
rect 79026 441922 79094 441978
rect 79150 441922 79218 441978
rect 79274 441922 79342 441978
rect 79398 441922 79494 441978
rect 78874 424350 79494 441922
rect 85168 436350 85488 436384
rect 85168 436294 85238 436350
rect 85294 436294 85362 436350
rect 85418 436294 85488 436350
rect 85168 436226 85488 436294
rect 85168 436170 85238 436226
rect 85294 436170 85362 436226
rect 85418 436170 85488 436226
rect 85168 436102 85488 436170
rect 85168 436046 85238 436102
rect 85294 436046 85362 436102
rect 85418 436046 85488 436102
rect 85168 435978 85488 436046
rect 85168 435922 85238 435978
rect 85294 435922 85362 435978
rect 85418 435922 85488 435978
rect 85168 435888 85488 435922
rect 93154 436350 93774 453922
rect 93154 436294 93250 436350
rect 93306 436294 93374 436350
rect 93430 436294 93498 436350
rect 93554 436294 93622 436350
rect 93678 436294 93774 436350
rect 93154 436226 93774 436294
rect 93154 436170 93250 436226
rect 93306 436170 93374 436226
rect 93430 436170 93498 436226
rect 93554 436170 93622 436226
rect 93678 436170 93774 436226
rect 93154 436102 93774 436170
rect 93154 436046 93250 436102
rect 93306 436046 93374 436102
rect 93430 436046 93498 436102
rect 93554 436046 93622 436102
rect 93678 436046 93774 436102
rect 93154 435978 93774 436046
rect 93154 435922 93250 435978
rect 93306 435922 93374 435978
rect 93430 435922 93498 435978
rect 93554 435922 93622 435978
rect 93678 435922 93774 435978
rect 78874 424294 78970 424350
rect 79026 424294 79094 424350
rect 79150 424294 79218 424350
rect 79274 424294 79342 424350
rect 79398 424294 79494 424350
rect 78874 424226 79494 424294
rect 78874 424170 78970 424226
rect 79026 424170 79094 424226
rect 79150 424170 79218 424226
rect 79274 424170 79342 424226
rect 79398 424170 79494 424226
rect 78874 424102 79494 424170
rect 78874 424046 78970 424102
rect 79026 424046 79094 424102
rect 79150 424046 79218 424102
rect 79274 424046 79342 424102
rect 79398 424046 79494 424102
rect 78874 423978 79494 424046
rect 78874 423922 78970 423978
rect 79026 423922 79094 423978
rect 79150 423922 79218 423978
rect 79274 423922 79342 423978
rect 79398 423922 79494 423978
rect 78874 406350 79494 423922
rect 85168 418350 85488 418384
rect 85168 418294 85238 418350
rect 85294 418294 85362 418350
rect 85418 418294 85488 418350
rect 85168 418226 85488 418294
rect 85168 418170 85238 418226
rect 85294 418170 85362 418226
rect 85418 418170 85488 418226
rect 85168 418102 85488 418170
rect 85168 418046 85238 418102
rect 85294 418046 85362 418102
rect 85418 418046 85488 418102
rect 85168 417978 85488 418046
rect 85168 417922 85238 417978
rect 85294 417922 85362 417978
rect 85418 417922 85488 417978
rect 85168 417888 85488 417922
rect 93154 418350 93774 435922
rect 93154 418294 93250 418350
rect 93306 418294 93374 418350
rect 93430 418294 93498 418350
rect 93554 418294 93622 418350
rect 93678 418294 93774 418350
rect 93154 418226 93774 418294
rect 93154 418170 93250 418226
rect 93306 418170 93374 418226
rect 93430 418170 93498 418226
rect 93554 418170 93622 418226
rect 93678 418170 93774 418226
rect 93154 418102 93774 418170
rect 93154 418046 93250 418102
rect 93306 418046 93374 418102
rect 93430 418046 93498 418102
rect 93554 418046 93622 418102
rect 93678 418046 93774 418102
rect 93154 417978 93774 418046
rect 93154 417922 93250 417978
rect 93306 417922 93374 417978
rect 93430 417922 93498 417978
rect 93554 417922 93622 417978
rect 93678 417922 93774 417978
rect 78874 406294 78970 406350
rect 79026 406294 79094 406350
rect 79150 406294 79218 406350
rect 79274 406294 79342 406350
rect 79398 406294 79494 406350
rect 78874 406226 79494 406294
rect 78874 406170 78970 406226
rect 79026 406170 79094 406226
rect 79150 406170 79218 406226
rect 79274 406170 79342 406226
rect 79398 406170 79494 406226
rect 78874 406102 79494 406170
rect 78874 406046 78970 406102
rect 79026 406046 79094 406102
rect 79150 406046 79218 406102
rect 79274 406046 79342 406102
rect 79398 406046 79494 406102
rect 78874 405978 79494 406046
rect 78874 405922 78970 405978
rect 79026 405922 79094 405978
rect 79150 405922 79218 405978
rect 79274 405922 79342 405978
rect 79398 405922 79494 405978
rect 78874 388350 79494 405922
rect 85168 400350 85488 400384
rect 85168 400294 85238 400350
rect 85294 400294 85362 400350
rect 85418 400294 85488 400350
rect 85168 400226 85488 400294
rect 85168 400170 85238 400226
rect 85294 400170 85362 400226
rect 85418 400170 85488 400226
rect 85168 400102 85488 400170
rect 85168 400046 85238 400102
rect 85294 400046 85362 400102
rect 85418 400046 85488 400102
rect 85168 399978 85488 400046
rect 85168 399922 85238 399978
rect 85294 399922 85362 399978
rect 85418 399922 85488 399978
rect 85168 399888 85488 399922
rect 93154 400350 93774 417922
rect 93154 400294 93250 400350
rect 93306 400294 93374 400350
rect 93430 400294 93498 400350
rect 93554 400294 93622 400350
rect 93678 400294 93774 400350
rect 93154 400226 93774 400294
rect 93154 400170 93250 400226
rect 93306 400170 93374 400226
rect 93430 400170 93498 400226
rect 93554 400170 93622 400226
rect 93678 400170 93774 400226
rect 93154 400102 93774 400170
rect 93154 400046 93250 400102
rect 93306 400046 93374 400102
rect 93430 400046 93498 400102
rect 93554 400046 93622 400102
rect 93678 400046 93774 400102
rect 93154 399978 93774 400046
rect 93154 399922 93250 399978
rect 93306 399922 93374 399978
rect 93430 399922 93498 399978
rect 93554 399922 93622 399978
rect 93678 399922 93774 399978
rect 78874 388294 78970 388350
rect 79026 388294 79094 388350
rect 79150 388294 79218 388350
rect 79274 388294 79342 388350
rect 79398 388294 79494 388350
rect 78874 388226 79494 388294
rect 78874 388170 78970 388226
rect 79026 388170 79094 388226
rect 79150 388170 79218 388226
rect 79274 388170 79342 388226
rect 79398 388170 79494 388226
rect 78874 388102 79494 388170
rect 78874 388046 78970 388102
rect 79026 388046 79094 388102
rect 79150 388046 79218 388102
rect 79274 388046 79342 388102
rect 79398 388046 79494 388102
rect 78874 387978 79494 388046
rect 78874 387922 78970 387978
rect 79026 387922 79094 387978
rect 79150 387922 79218 387978
rect 79274 387922 79342 387978
rect 79398 387922 79494 387978
rect 78874 370350 79494 387922
rect 85168 382350 85488 382384
rect 85168 382294 85238 382350
rect 85294 382294 85362 382350
rect 85418 382294 85488 382350
rect 85168 382226 85488 382294
rect 85168 382170 85238 382226
rect 85294 382170 85362 382226
rect 85418 382170 85488 382226
rect 85168 382102 85488 382170
rect 85168 382046 85238 382102
rect 85294 382046 85362 382102
rect 85418 382046 85488 382102
rect 85168 381978 85488 382046
rect 85168 381922 85238 381978
rect 85294 381922 85362 381978
rect 85418 381922 85488 381978
rect 85168 381888 85488 381922
rect 93154 382350 93774 399922
rect 93154 382294 93250 382350
rect 93306 382294 93374 382350
rect 93430 382294 93498 382350
rect 93554 382294 93622 382350
rect 93678 382294 93774 382350
rect 93154 382226 93774 382294
rect 93154 382170 93250 382226
rect 93306 382170 93374 382226
rect 93430 382170 93498 382226
rect 93554 382170 93622 382226
rect 93678 382170 93774 382226
rect 93154 382102 93774 382170
rect 93154 382046 93250 382102
rect 93306 382046 93374 382102
rect 93430 382046 93498 382102
rect 93554 382046 93622 382102
rect 93678 382046 93774 382102
rect 93154 381978 93774 382046
rect 93154 381922 93250 381978
rect 93306 381922 93374 381978
rect 93430 381922 93498 381978
rect 93554 381922 93622 381978
rect 93678 381922 93774 381978
rect 78874 370294 78970 370350
rect 79026 370294 79094 370350
rect 79150 370294 79218 370350
rect 79274 370294 79342 370350
rect 79398 370294 79494 370350
rect 78874 370226 79494 370294
rect 78874 370170 78970 370226
rect 79026 370170 79094 370226
rect 79150 370170 79218 370226
rect 79274 370170 79342 370226
rect 79398 370170 79494 370226
rect 78874 370102 79494 370170
rect 78874 370046 78970 370102
rect 79026 370046 79094 370102
rect 79150 370046 79218 370102
rect 79274 370046 79342 370102
rect 79398 370046 79494 370102
rect 78874 369978 79494 370046
rect 78874 369922 78970 369978
rect 79026 369922 79094 369978
rect 79150 369922 79218 369978
rect 79274 369922 79342 369978
rect 79398 369922 79494 369978
rect 78874 352350 79494 369922
rect 85168 364350 85488 364384
rect 85168 364294 85238 364350
rect 85294 364294 85362 364350
rect 85418 364294 85488 364350
rect 85168 364226 85488 364294
rect 85168 364170 85238 364226
rect 85294 364170 85362 364226
rect 85418 364170 85488 364226
rect 85168 364102 85488 364170
rect 85168 364046 85238 364102
rect 85294 364046 85362 364102
rect 85418 364046 85488 364102
rect 85168 363978 85488 364046
rect 85168 363922 85238 363978
rect 85294 363922 85362 363978
rect 85418 363922 85488 363978
rect 85168 363888 85488 363922
rect 93154 364350 93774 381922
rect 93154 364294 93250 364350
rect 93306 364294 93374 364350
rect 93430 364294 93498 364350
rect 93554 364294 93622 364350
rect 93678 364294 93774 364350
rect 93154 364226 93774 364294
rect 93154 364170 93250 364226
rect 93306 364170 93374 364226
rect 93430 364170 93498 364226
rect 93554 364170 93622 364226
rect 93678 364170 93774 364226
rect 93154 364102 93774 364170
rect 93154 364046 93250 364102
rect 93306 364046 93374 364102
rect 93430 364046 93498 364102
rect 93554 364046 93622 364102
rect 93678 364046 93774 364102
rect 93154 363978 93774 364046
rect 93154 363922 93250 363978
rect 93306 363922 93374 363978
rect 93430 363922 93498 363978
rect 93554 363922 93622 363978
rect 93678 363922 93774 363978
rect 78874 352294 78970 352350
rect 79026 352294 79094 352350
rect 79150 352294 79218 352350
rect 79274 352294 79342 352350
rect 79398 352294 79494 352350
rect 78874 352226 79494 352294
rect 78874 352170 78970 352226
rect 79026 352170 79094 352226
rect 79150 352170 79218 352226
rect 79274 352170 79342 352226
rect 79398 352170 79494 352226
rect 78874 352102 79494 352170
rect 78874 352046 78970 352102
rect 79026 352046 79094 352102
rect 79150 352046 79218 352102
rect 79274 352046 79342 352102
rect 79398 352046 79494 352102
rect 78874 351978 79494 352046
rect 78874 351922 78970 351978
rect 79026 351922 79094 351978
rect 79150 351922 79218 351978
rect 79274 351922 79342 351978
rect 79398 351922 79494 351978
rect 78874 334350 79494 351922
rect 85168 346350 85488 346384
rect 85168 346294 85238 346350
rect 85294 346294 85362 346350
rect 85418 346294 85488 346350
rect 85168 346226 85488 346294
rect 85168 346170 85238 346226
rect 85294 346170 85362 346226
rect 85418 346170 85488 346226
rect 85168 346102 85488 346170
rect 85168 346046 85238 346102
rect 85294 346046 85362 346102
rect 85418 346046 85488 346102
rect 85168 345978 85488 346046
rect 85168 345922 85238 345978
rect 85294 345922 85362 345978
rect 85418 345922 85488 345978
rect 85168 345888 85488 345922
rect 93154 346350 93774 363922
rect 93154 346294 93250 346350
rect 93306 346294 93374 346350
rect 93430 346294 93498 346350
rect 93554 346294 93622 346350
rect 93678 346294 93774 346350
rect 93154 346226 93774 346294
rect 93154 346170 93250 346226
rect 93306 346170 93374 346226
rect 93430 346170 93498 346226
rect 93554 346170 93622 346226
rect 93678 346170 93774 346226
rect 93154 346102 93774 346170
rect 93154 346046 93250 346102
rect 93306 346046 93374 346102
rect 93430 346046 93498 346102
rect 93554 346046 93622 346102
rect 93678 346046 93774 346102
rect 93154 345978 93774 346046
rect 93154 345922 93250 345978
rect 93306 345922 93374 345978
rect 93430 345922 93498 345978
rect 93554 345922 93622 345978
rect 93678 345922 93774 345978
rect 78874 334294 78970 334350
rect 79026 334294 79094 334350
rect 79150 334294 79218 334350
rect 79274 334294 79342 334350
rect 79398 334294 79494 334350
rect 78874 334226 79494 334294
rect 78874 334170 78970 334226
rect 79026 334170 79094 334226
rect 79150 334170 79218 334226
rect 79274 334170 79342 334226
rect 79398 334170 79494 334226
rect 78874 334102 79494 334170
rect 78874 334046 78970 334102
rect 79026 334046 79094 334102
rect 79150 334046 79218 334102
rect 79274 334046 79342 334102
rect 79398 334046 79494 334102
rect 78874 333978 79494 334046
rect 78874 333922 78970 333978
rect 79026 333922 79094 333978
rect 79150 333922 79218 333978
rect 79274 333922 79342 333978
rect 79398 333922 79494 333978
rect 78874 316350 79494 333922
rect 85168 328350 85488 328384
rect 85168 328294 85238 328350
rect 85294 328294 85362 328350
rect 85418 328294 85488 328350
rect 85168 328226 85488 328294
rect 85168 328170 85238 328226
rect 85294 328170 85362 328226
rect 85418 328170 85488 328226
rect 85168 328102 85488 328170
rect 85168 328046 85238 328102
rect 85294 328046 85362 328102
rect 85418 328046 85488 328102
rect 85168 327978 85488 328046
rect 85168 327922 85238 327978
rect 85294 327922 85362 327978
rect 85418 327922 85488 327978
rect 85168 327888 85488 327922
rect 93154 328350 93774 345922
rect 93154 328294 93250 328350
rect 93306 328294 93374 328350
rect 93430 328294 93498 328350
rect 93554 328294 93622 328350
rect 93678 328294 93774 328350
rect 93154 328226 93774 328294
rect 93154 328170 93250 328226
rect 93306 328170 93374 328226
rect 93430 328170 93498 328226
rect 93554 328170 93622 328226
rect 93678 328170 93774 328226
rect 93154 328102 93774 328170
rect 93154 328046 93250 328102
rect 93306 328046 93374 328102
rect 93430 328046 93498 328102
rect 93554 328046 93622 328102
rect 93678 328046 93774 328102
rect 93154 327978 93774 328046
rect 93154 327922 93250 327978
rect 93306 327922 93374 327978
rect 93430 327922 93498 327978
rect 93554 327922 93622 327978
rect 93678 327922 93774 327978
rect 78874 316294 78970 316350
rect 79026 316294 79094 316350
rect 79150 316294 79218 316350
rect 79274 316294 79342 316350
rect 79398 316294 79494 316350
rect 78874 316226 79494 316294
rect 78874 316170 78970 316226
rect 79026 316170 79094 316226
rect 79150 316170 79218 316226
rect 79274 316170 79342 316226
rect 79398 316170 79494 316226
rect 78874 316102 79494 316170
rect 78874 316046 78970 316102
rect 79026 316046 79094 316102
rect 79150 316046 79218 316102
rect 79274 316046 79342 316102
rect 79398 316046 79494 316102
rect 78874 315978 79494 316046
rect 78874 315922 78970 315978
rect 79026 315922 79094 315978
rect 79150 315922 79218 315978
rect 79274 315922 79342 315978
rect 79398 315922 79494 315978
rect 78874 298350 79494 315922
rect 85168 310350 85488 310384
rect 85168 310294 85238 310350
rect 85294 310294 85362 310350
rect 85418 310294 85488 310350
rect 85168 310226 85488 310294
rect 85168 310170 85238 310226
rect 85294 310170 85362 310226
rect 85418 310170 85488 310226
rect 85168 310102 85488 310170
rect 85168 310046 85238 310102
rect 85294 310046 85362 310102
rect 85418 310046 85488 310102
rect 85168 309978 85488 310046
rect 85168 309922 85238 309978
rect 85294 309922 85362 309978
rect 85418 309922 85488 309978
rect 85168 309888 85488 309922
rect 93154 310350 93774 327922
rect 93154 310294 93250 310350
rect 93306 310294 93374 310350
rect 93430 310294 93498 310350
rect 93554 310294 93622 310350
rect 93678 310294 93774 310350
rect 93154 310226 93774 310294
rect 93154 310170 93250 310226
rect 93306 310170 93374 310226
rect 93430 310170 93498 310226
rect 93554 310170 93622 310226
rect 93678 310170 93774 310226
rect 93154 310102 93774 310170
rect 93154 310046 93250 310102
rect 93306 310046 93374 310102
rect 93430 310046 93498 310102
rect 93554 310046 93622 310102
rect 93678 310046 93774 310102
rect 93154 309978 93774 310046
rect 93154 309922 93250 309978
rect 93306 309922 93374 309978
rect 93430 309922 93498 309978
rect 93554 309922 93622 309978
rect 93678 309922 93774 309978
rect 78874 298294 78970 298350
rect 79026 298294 79094 298350
rect 79150 298294 79218 298350
rect 79274 298294 79342 298350
rect 79398 298294 79494 298350
rect 78874 298226 79494 298294
rect 78874 298170 78970 298226
rect 79026 298170 79094 298226
rect 79150 298170 79218 298226
rect 79274 298170 79342 298226
rect 79398 298170 79494 298226
rect 78874 298102 79494 298170
rect 78874 298046 78970 298102
rect 79026 298046 79094 298102
rect 79150 298046 79218 298102
rect 79274 298046 79342 298102
rect 79398 298046 79494 298102
rect 78874 297978 79494 298046
rect 78874 297922 78970 297978
rect 79026 297922 79094 297978
rect 79150 297922 79218 297978
rect 79274 297922 79342 297978
rect 79398 297922 79494 297978
rect 78874 280350 79494 297922
rect 85168 292350 85488 292384
rect 85168 292294 85238 292350
rect 85294 292294 85362 292350
rect 85418 292294 85488 292350
rect 85168 292226 85488 292294
rect 85168 292170 85238 292226
rect 85294 292170 85362 292226
rect 85418 292170 85488 292226
rect 85168 292102 85488 292170
rect 85168 292046 85238 292102
rect 85294 292046 85362 292102
rect 85418 292046 85488 292102
rect 85168 291978 85488 292046
rect 85168 291922 85238 291978
rect 85294 291922 85362 291978
rect 85418 291922 85488 291978
rect 85168 291888 85488 291922
rect 93154 292350 93774 309922
rect 93154 292294 93250 292350
rect 93306 292294 93374 292350
rect 93430 292294 93498 292350
rect 93554 292294 93622 292350
rect 93678 292294 93774 292350
rect 93154 292226 93774 292294
rect 93154 292170 93250 292226
rect 93306 292170 93374 292226
rect 93430 292170 93498 292226
rect 93554 292170 93622 292226
rect 93678 292170 93774 292226
rect 93154 292102 93774 292170
rect 93154 292046 93250 292102
rect 93306 292046 93374 292102
rect 93430 292046 93498 292102
rect 93554 292046 93622 292102
rect 93678 292046 93774 292102
rect 93154 291978 93774 292046
rect 93154 291922 93250 291978
rect 93306 291922 93374 291978
rect 93430 291922 93498 291978
rect 93554 291922 93622 291978
rect 93678 291922 93774 291978
rect 78874 280294 78970 280350
rect 79026 280294 79094 280350
rect 79150 280294 79218 280350
rect 79274 280294 79342 280350
rect 79398 280294 79494 280350
rect 78874 280226 79494 280294
rect 78874 280170 78970 280226
rect 79026 280170 79094 280226
rect 79150 280170 79218 280226
rect 79274 280170 79342 280226
rect 79398 280170 79494 280226
rect 78874 280102 79494 280170
rect 78874 280046 78970 280102
rect 79026 280046 79094 280102
rect 79150 280046 79218 280102
rect 79274 280046 79342 280102
rect 79398 280046 79494 280102
rect 78874 279978 79494 280046
rect 78874 279922 78970 279978
rect 79026 279922 79094 279978
rect 79150 279922 79218 279978
rect 79274 279922 79342 279978
rect 79398 279922 79494 279978
rect 78874 262350 79494 279922
rect 85168 274350 85488 274384
rect 85168 274294 85238 274350
rect 85294 274294 85362 274350
rect 85418 274294 85488 274350
rect 85168 274226 85488 274294
rect 85168 274170 85238 274226
rect 85294 274170 85362 274226
rect 85418 274170 85488 274226
rect 85168 274102 85488 274170
rect 85168 274046 85238 274102
rect 85294 274046 85362 274102
rect 85418 274046 85488 274102
rect 85168 273978 85488 274046
rect 85168 273922 85238 273978
rect 85294 273922 85362 273978
rect 85418 273922 85488 273978
rect 85168 273888 85488 273922
rect 93154 274350 93774 291922
rect 93154 274294 93250 274350
rect 93306 274294 93374 274350
rect 93430 274294 93498 274350
rect 93554 274294 93622 274350
rect 93678 274294 93774 274350
rect 93154 274226 93774 274294
rect 93154 274170 93250 274226
rect 93306 274170 93374 274226
rect 93430 274170 93498 274226
rect 93554 274170 93622 274226
rect 93678 274170 93774 274226
rect 93154 274102 93774 274170
rect 93154 274046 93250 274102
rect 93306 274046 93374 274102
rect 93430 274046 93498 274102
rect 93554 274046 93622 274102
rect 93678 274046 93774 274102
rect 93154 273978 93774 274046
rect 93154 273922 93250 273978
rect 93306 273922 93374 273978
rect 93430 273922 93498 273978
rect 93554 273922 93622 273978
rect 93678 273922 93774 273978
rect 78874 262294 78970 262350
rect 79026 262294 79094 262350
rect 79150 262294 79218 262350
rect 79274 262294 79342 262350
rect 79398 262294 79494 262350
rect 78874 262226 79494 262294
rect 78874 262170 78970 262226
rect 79026 262170 79094 262226
rect 79150 262170 79218 262226
rect 79274 262170 79342 262226
rect 79398 262170 79494 262226
rect 78874 262102 79494 262170
rect 78874 262046 78970 262102
rect 79026 262046 79094 262102
rect 79150 262046 79218 262102
rect 79274 262046 79342 262102
rect 79398 262046 79494 262102
rect 78874 261978 79494 262046
rect 78874 261922 78970 261978
rect 79026 261922 79094 261978
rect 79150 261922 79218 261978
rect 79274 261922 79342 261978
rect 79398 261922 79494 261978
rect 78874 244350 79494 261922
rect 85168 256350 85488 256384
rect 85168 256294 85238 256350
rect 85294 256294 85362 256350
rect 85418 256294 85488 256350
rect 85168 256226 85488 256294
rect 85168 256170 85238 256226
rect 85294 256170 85362 256226
rect 85418 256170 85488 256226
rect 85168 256102 85488 256170
rect 85168 256046 85238 256102
rect 85294 256046 85362 256102
rect 85418 256046 85488 256102
rect 85168 255978 85488 256046
rect 85168 255922 85238 255978
rect 85294 255922 85362 255978
rect 85418 255922 85488 255978
rect 85168 255888 85488 255922
rect 93154 256350 93774 273922
rect 93154 256294 93250 256350
rect 93306 256294 93374 256350
rect 93430 256294 93498 256350
rect 93554 256294 93622 256350
rect 93678 256294 93774 256350
rect 93154 256226 93774 256294
rect 93154 256170 93250 256226
rect 93306 256170 93374 256226
rect 93430 256170 93498 256226
rect 93554 256170 93622 256226
rect 93678 256170 93774 256226
rect 93154 256102 93774 256170
rect 93154 256046 93250 256102
rect 93306 256046 93374 256102
rect 93430 256046 93498 256102
rect 93554 256046 93622 256102
rect 93678 256046 93774 256102
rect 93154 255978 93774 256046
rect 93154 255922 93250 255978
rect 93306 255922 93374 255978
rect 93430 255922 93498 255978
rect 93554 255922 93622 255978
rect 93678 255922 93774 255978
rect 78874 244294 78970 244350
rect 79026 244294 79094 244350
rect 79150 244294 79218 244350
rect 79274 244294 79342 244350
rect 79398 244294 79494 244350
rect 78874 244226 79494 244294
rect 78874 244170 78970 244226
rect 79026 244170 79094 244226
rect 79150 244170 79218 244226
rect 79274 244170 79342 244226
rect 79398 244170 79494 244226
rect 78874 244102 79494 244170
rect 78874 244046 78970 244102
rect 79026 244046 79094 244102
rect 79150 244046 79218 244102
rect 79274 244046 79342 244102
rect 79398 244046 79494 244102
rect 78874 243978 79494 244046
rect 78874 243922 78970 243978
rect 79026 243922 79094 243978
rect 79150 243922 79218 243978
rect 79274 243922 79342 243978
rect 79398 243922 79494 243978
rect 78874 226350 79494 243922
rect 85168 238350 85488 238384
rect 85168 238294 85238 238350
rect 85294 238294 85362 238350
rect 85418 238294 85488 238350
rect 85168 238226 85488 238294
rect 85168 238170 85238 238226
rect 85294 238170 85362 238226
rect 85418 238170 85488 238226
rect 85168 238102 85488 238170
rect 85168 238046 85238 238102
rect 85294 238046 85362 238102
rect 85418 238046 85488 238102
rect 85168 237978 85488 238046
rect 85168 237922 85238 237978
rect 85294 237922 85362 237978
rect 85418 237922 85488 237978
rect 85168 237888 85488 237922
rect 93154 238350 93774 255922
rect 93154 238294 93250 238350
rect 93306 238294 93374 238350
rect 93430 238294 93498 238350
rect 93554 238294 93622 238350
rect 93678 238294 93774 238350
rect 93154 238226 93774 238294
rect 93154 238170 93250 238226
rect 93306 238170 93374 238226
rect 93430 238170 93498 238226
rect 93554 238170 93622 238226
rect 93678 238170 93774 238226
rect 93154 238102 93774 238170
rect 93154 238046 93250 238102
rect 93306 238046 93374 238102
rect 93430 238046 93498 238102
rect 93554 238046 93622 238102
rect 93678 238046 93774 238102
rect 93154 237978 93774 238046
rect 93154 237922 93250 237978
rect 93306 237922 93374 237978
rect 93430 237922 93498 237978
rect 93554 237922 93622 237978
rect 93678 237922 93774 237978
rect 78874 226294 78970 226350
rect 79026 226294 79094 226350
rect 79150 226294 79218 226350
rect 79274 226294 79342 226350
rect 79398 226294 79494 226350
rect 78874 226226 79494 226294
rect 78874 226170 78970 226226
rect 79026 226170 79094 226226
rect 79150 226170 79218 226226
rect 79274 226170 79342 226226
rect 79398 226170 79494 226226
rect 78874 226102 79494 226170
rect 78874 226046 78970 226102
rect 79026 226046 79094 226102
rect 79150 226046 79218 226102
rect 79274 226046 79342 226102
rect 79398 226046 79494 226102
rect 78874 225978 79494 226046
rect 78874 225922 78970 225978
rect 79026 225922 79094 225978
rect 79150 225922 79218 225978
rect 79274 225922 79342 225978
rect 79398 225922 79494 225978
rect 78874 208350 79494 225922
rect 85168 220350 85488 220384
rect 85168 220294 85238 220350
rect 85294 220294 85362 220350
rect 85418 220294 85488 220350
rect 85168 220226 85488 220294
rect 85168 220170 85238 220226
rect 85294 220170 85362 220226
rect 85418 220170 85488 220226
rect 85168 220102 85488 220170
rect 85168 220046 85238 220102
rect 85294 220046 85362 220102
rect 85418 220046 85488 220102
rect 85168 219978 85488 220046
rect 85168 219922 85238 219978
rect 85294 219922 85362 219978
rect 85418 219922 85488 219978
rect 85168 219888 85488 219922
rect 93154 220350 93774 237922
rect 93154 220294 93250 220350
rect 93306 220294 93374 220350
rect 93430 220294 93498 220350
rect 93554 220294 93622 220350
rect 93678 220294 93774 220350
rect 93154 220226 93774 220294
rect 93154 220170 93250 220226
rect 93306 220170 93374 220226
rect 93430 220170 93498 220226
rect 93554 220170 93622 220226
rect 93678 220170 93774 220226
rect 93154 220102 93774 220170
rect 93154 220046 93250 220102
rect 93306 220046 93374 220102
rect 93430 220046 93498 220102
rect 93554 220046 93622 220102
rect 93678 220046 93774 220102
rect 93154 219978 93774 220046
rect 93154 219922 93250 219978
rect 93306 219922 93374 219978
rect 93430 219922 93498 219978
rect 93554 219922 93622 219978
rect 93678 219922 93774 219978
rect 78874 208294 78970 208350
rect 79026 208294 79094 208350
rect 79150 208294 79218 208350
rect 79274 208294 79342 208350
rect 79398 208294 79494 208350
rect 78874 208226 79494 208294
rect 78874 208170 78970 208226
rect 79026 208170 79094 208226
rect 79150 208170 79218 208226
rect 79274 208170 79342 208226
rect 79398 208170 79494 208226
rect 78874 208102 79494 208170
rect 78874 208046 78970 208102
rect 79026 208046 79094 208102
rect 79150 208046 79218 208102
rect 79274 208046 79342 208102
rect 79398 208046 79494 208102
rect 78874 207978 79494 208046
rect 78874 207922 78970 207978
rect 79026 207922 79094 207978
rect 79150 207922 79218 207978
rect 79274 207922 79342 207978
rect 79398 207922 79494 207978
rect 78874 190350 79494 207922
rect 85168 202350 85488 202384
rect 85168 202294 85238 202350
rect 85294 202294 85362 202350
rect 85418 202294 85488 202350
rect 85168 202226 85488 202294
rect 85168 202170 85238 202226
rect 85294 202170 85362 202226
rect 85418 202170 85488 202226
rect 85168 202102 85488 202170
rect 85168 202046 85238 202102
rect 85294 202046 85362 202102
rect 85418 202046 85488 202102
rect 85168 201978 85488 202046
rect 85168 201922 85238 201978
rect 85294 201922 85362 201978
rect 85418 201922 85488 201978
rect 85168 201888 85488 201922
rect 93154 202350 93774 219922
rect 93154 202294 93250 202350
rect 93306 202294 93374 202350
rect 93430 202294 93498 202350
rect 93554 202294 93622 202350
rect 93678 202294 93774 202350
rect 93154 202226 93774 202294
rect 93154 202170 93250 202226
rect 93306 202170 93374 202226
rect 93430 202170 93498 202226
rect 93554 202170 93622 202226
rect 93678 202170 93774 202226
rect 93154 202102 93774 202170
rect 93154 202046 93250 202102
rect 93306 202046 93374 202102
rect 93430 202046 93498 202102
rect 93554 202046 93622 202102
rect 93678 202046 93774 202102
rect 93154 201978 93774 202046
rect 93154 201922 93250 201978
rect 93306 201922 93374 201978
rect 93430 201922 93498 201978
rect 93554 201922 93622 201978
rect 93678 201922 93774 201978
rect 78874 190294 78970 190350
rect 79026 190294 79094 190350
rect 79150 190294 79218 190350
rect 79274 190294 79342 190350
rect 79398 190294 79494 190350
rect 78874 190226 79494 190294
rect 78874 190170 78970 190226
rect 79026 190170 79094 190226
rect 79150 190170 79218 190226
rect 79274 190170 79342 190226
rect 79398 190170 79494 190226
rect 78874 190102 79494 190170
rect 78874 190046 78970 190102
rect 79026 190046 79094 190102
rect 79150 190046 79218 190102
rect 79274 190046 79342 190102
rect 79398 190046 79494 190102
rect 78874 189978 79494 190046
rect 78874 189922 78970 189978
rect 79026 189922 79094 189978
rect 79150 189922 79218 189978
rect 79274 189922 79342 189978
rect 79398 189922 79494 189978
rect 78874 172350 79494 189922
rect 85168 184350 85488 184384
rect 85168 184294 85238 184350
rect 85294 184294 85362 184350
rect 85418 184294 85488 184350
rect 85168 184226 85488 184294
rect 85168 184170 85238 184226
rect 85294 184170 85362 184226
rect 85418 184170 85488 184226
rect 85168 184102 85488 184170
rect 85168 184046 85238 184102
rect 85294 184046 85362 184102
rect 85418 184046 85488 184102
rect 85168 183978 85488 184046
rect 85168 183922 85238 183978
rect 85294 183922 85362 183978
rect 85418 183922 85488 183978
rect 85168 183888 85488 183922
rect 93154 184350 93774 201922
rect 93154 184294 93250 184350
rect 93306 184294 93374 184350
rect 93430 184294 93498 184350
rect 93554 184294 93622 184350
rect 93678 184294 93774 184350
rect 93154 184226 93774 184294
rect 93154 184170 93250 184226
rect 93306 184170 93374 184226
rect 93430 184170 93498 184226
rect 93554 184170 93622 184226
rect 93678 184170 93774 184226
rect 93154 184102 93774 184170
rect 93154 184046 93250 184102
rect 93306 184046 93374 184102
rect 93430 184046 93498 184102
rect 93554 184046 93622 184102
rect 93678 184046 93774 184102
rect 93154 183978 93774 184046
rect 93154 183922 93250 183978
rect 93306 183922 93374 183978
rect 93430 183922 93498 183978
rect 93554 183922 93622 183978
rect 93678 183922 93774 183978
rect 78874 172294 78970 172350
rect 79026 172294 79094 172350
rect 79150 172294 79218 172350
rect 79274 172294 79342 172350
rect 79398 172294 79494 172350
rect 78874 172226 79494 172294
rect 78874 172170 78970 172226
rect 79026 172170 79094 172226
rect 79150 172170 79218 172226
rect 79274 172170 79342 172226
rect 79398 172170 79494 172226
rect 78874 172102 79494 172170
rect 78874 172046 78970 172102
rect 79026 172046 79094 172102
rect 79150 172046 79218 172102
rect 79274 172046 79342 172102
rect 79398 172046 79494 172102
rect 78874 171978 79494 172046
rect 78874 171922 78970 171978
rect 79026 171922 79094 171978
rect 79150 171922 79218 171978
rect 79274 171922 79342 171978
rect 79398 171922 79494 171978
rect 78874 154350 79494 171922
rect 85168 166350 85488 166384
rect 85168 166294 85238 166350
rect 85294 166294 85362 166350
rect 85418 166294 85488 166350
rect 85168 166226 85488 166294
rect 85168 166170 85238 166226
rect 85294 166170 85362 166226
rect 85418 166170 85488 166226
rect 85168 166102 85488 166170
rect 85168 166046 85238 166102
rect 85294 166046 85362 166102
rect 85418 166046 85488 166102
rect 85168 165978 85488 166046
rect 85168 165922 85238 165978
rect 85294 165922 85362 165978
rect 85418 165922 85488 165978
rect 85168 165888 85488 165922
rect 93154 166350 93774 183922
rect 93154 166294 93250 166350
rect 93306 166294 93374 166350
rect 93430 166294 93498 166350
rect 93554 166294 93622 166350
rect 93678 166294 93774 166350
rect 93154 166226 93774 166294
rect 93154 166170 93250 166226
rect 93306 166170 93374 166226
rect 93430 166170 93498 166226
rect 93554 166170 93622 166226
rect 93678 166170 93774 166226
rect 93154 166102 93774 166170
rect 93154 166046 93250 166102
rect 93306 166046 93374 166102
rect 93430 166046 93498 166102
rect 93554 166046 93622 166102
rect 93678 166046 93774 166102
rect 93154 165978 93774 166046
rect 93154 165922 93250 165978
rect 93306 165922 93374 165978
rect 93430 165922 93498 165978
rect 93554 165922 93622 165978
rect 93678 165922 93774 165978
rect 78874 154294 78970 154350
rect 79026 154294 79094 154350
rect 79150 154294 79218 154350
rect 79274 154294 79342 154350
rect 79398 154294 79494 154350
rect 78874 154226 79494 154294
rect 78874 154170 78970 154226
rect 79026 154170 79094 154226
rect 79150 154170 79218 154226
rect 79274 154170 79342 154226
rect 79398 154170 79494 154226
rect 78874 154102 79494 154170
rect 78874 154046 78970 154102
rect 79026 154046 79094 154102
rect 79150 154046 79218 154102
rect 79274 154046 79342 154102
rect 79398 154046 79494 154102
rect 78874 153978 79494 154046
rect 78874 153922 78970 153978
rect 79026 153922 79094 153978
rect 79150 153922 79218 153978
rect 79274 153922 79342 153978
rect 79398 153922 79494 153978
rect 78874 136350 79494 153922
rect 85168 148350 85488 148384
rect 85168 148294 85238 148350
rect 85294 148294 85362 148350
rect 85418 148294 85488 148350
rect 85168 148226 85488 148294
rect 85168 148170 85238 148226
rect 85294 148170 85362 148226
rect 85418 148170 85488 148226
rect 85168 148102 85488 148170
rect 85168 148046 85238 148102
rect 85294 148046 85362 148102
rect 85418 148046 85488 148102
rect 85168 147978 85488 148046
rect 85168 147922 85238 147978
rect 85294 147922 85362 147978
rect 85418 147922 85488 147978
rect 85168 147888 85488 147922
rect 93154 148350 93774 165922
rect 93154 148294 93250 148350
rect 93306 148294 93374 148350
rect 93430 148294 93498 148350
rect 93554 148294 93622 148350
rect 93678 148294 93774 148350
rect 93154 148226 93774 148294
rect 93154 148170 93250 148226
rect 93306 148170 93374 148226
rect 93430 148170 93498 148226
rect 93554 148170 93622 148226
rect 93678 148170 93774 148226
rect 93154 148102 93774 148170
rect 93154 148046 93250 148102
rect 93306 148046 93374 148102
rect 93430 148046 93498 148102
rect 93554 148046 93622 148102
rect 93678 148046 93774 148102
rect 93154 147978 93774 148046
rect 93154 147922 93250 147978
rect 93306 147922 93374 147978
rect 93430 147922 93498 147978
rect 93554 147922 93622 147978
rect 93678 147922 93774 147978
rect 78874 136294 78970 136350
rect 79026 136294 79094 136350
rect 79150 136294 79218 136350
rect 79274 136294 79342 136350
rect 79398 136294 79494 136350
rect 78874 136226 79494 136294
rect 78874 136170 78970 136226
rect 79026 136170 79094 136226
rect 79150 136170 79218 136226
rect 79274 136170 79342 136226
rect 79398 136170 79494 136226
rect 78874 136102 79494 136170
rect 78874 136046 78970 136102
rect 79026 136046 79094 136102
rect 79150 136046 79218 136102
rect 79274 136046 79342 136102
rect 79398 136046 79494 136102
rect 78874 135978 79494 136046
rect 78874 135922 78970 135978
rect 79026 135922 79094 135978
rect 79150 135922 79218 135978
rect 79274 135922 79342 135978
rect 79398 135922 79494 135978
rect 78874 118350 79494 135922
rect 85168 130350 85488 130384
rect 85168 130294 85238 130350
rect 85294 130294 85362 130350
rect 85418 130294 85488 130350
rect 85168 130226 85488 130294
rect 85168 130170 85238 130226
rect 85294 130170 85362 130226
rect 85418 130170 85488 130226
rect 85168 130102 85488 130170
rect 85168 130046 85238 130102
rect 85294 130046 85362 130102
rect 85418 130046 85488 130102
rect 85168 129978 85488 130046
rect 85168 129922 85238 129978
rect 85294 129922 85362 129978
rect 85418 129922 85488 129978
rect 85168 129888 85488 129922
rect 93154 130350 93774 147922
rect 93154 130294 93250 130350
rect 93306 130294 93374 130350
rect 93430 130294 93498 130350
rect 93554 130294 93622 130350
rect 93678 130294 93774 130350
rect 93154 130226 93774 130294
rect 93154 130170 93250 130226
rect 93306 130170 93374 130226
rect 93430 130170 93498 130226
rect 93554 130170 93622 130226
rect 93678 130170 93774 130226
rect 93154 130102 93774 130170
rect 93154 130046 93250 130102
rect 93306 130046 93374 130102
rect 93430 130046 93498 130102
rect 93554 130046 93622 130102
rect 93678 130046 93774 130102
rect 93154 129978 93774 130046
rect 93154 129922 93250 129978
rect 93306 129922 93374 129978
rect 93430 129922 93498 129978
rect 93554 129922 93622 129978
rect 93678 129922 93774 129978
rect 78874 118294 78970 118350
rect 79026 118294 79094 118350
rect 79150 118294 79218 118350
rect 79274 118294 79342 118350
rect 79398 118294 79494 118350
rect 78874 118226 79494 118294
rect 78874 118170 78970 118226
rect 79026 118170 79094 118226
rect 79150 118170 79218 118226
rect 79274 118170 79342 118226
rect 79398 118170 79494 118226
rect 78874 118102 79494 118170
rect 78874 118046 78970 118102
rect 79026 118046 79094 118102
rect 79150 118046 79218 118102
rect 79274 118046 79342 118102
rect 79398 118046 79494 118102
rect 78874 117978 79494 118046
rect 78874 117922 78970 117978
rect 79026 117922 79094 117978
rect 79150 117922 79218 117978
rect 79274 117922 79342 117978
rect 79398 117922 79494 117978
rect 78874 100350 79494 117922
rect 85168 112350 85488 112384
rect 85168 112294 85238 112350
rect 85294 112294 85362 112350
rect 85418 112294 85488 112350
rect 85168 112226 85488 112294
rect 85168 112170 85238 112226
rect 85294 112170 85362 112226
rect 85418 112170 85488 112226
rect 85168 112102 85488 112170
rect 85168 112046 85238 112102
rect 85294 112046 85362 112102
rect 85418 112046 85488 112102
rect 85168 111978 85488 112046
rect 85168 111922 85238 111978
rect 85294 111922 85362 111978
rect 85418 111922 85488 111978
rect 85168 111888 85488 111922
rect 93154 112350 93774 129922
rect 93154 112294 93250 112350
rect 93306 112294 93374 112350
rect 93430 112294 93498 112350
rect 93554 112294 93622 112350
rect 93678 112294 93774 112350
rect 93154 112226 93774 112294
rect 93154 112170 93250 112226
rect 93306 112170 93374 112226
rect 93430 112170 93498 112226
rect 93554 112170 93622 112226
rect 93678 112170 93774 112226
rect 93154 112102 93774 112170
rect 93154 112046 93250 112102
rect 93306 112046 93374 112102
rect 93430 112046 93498 112102
rect 93554 112046 93622 112102
rect 93678 112046 93774 112102
rect 93154 111978 93774 112046
rect 93154 111922 93250 111978
rect 93306 111922 93374 111978
rect 93430 111922 93498 111978
rect 93554 111922 93622 111978
rect 93678 111922 93774 111978
rect 78874 100294 78970 100350
rect 79026 100294 79094 100350
rect 79150 100294 79218 100350
rect 79274 100294 79342 100350
rect 79398 100294 79494 100350
rect 78874 100226 79494 100294
rect 78874 100170 78970 100226
rect 79026 100170 79094 100226
rect 79150 100170 79218 100226
rect 79274 100170 79342 100226
rect 79398 100170 79494 100226
rect 78874 100102 79494 100170
rect 78874 100046 78970 100102
rect 79026 100046 79094 100102
rect 79150 100046 79218 100102
rect 79274 100046 79342 100102
rect 79398 100046 79494 100102
rect 78874 99978 79494 100046
rect 78874 99922 78970 99978
rect 79026 99922 79094 99978
rect 79150 99922 79218 99978
rect 79274 99922 79342 99978
rect 79398 99922 79494 99978
rect 78874 82350 79494 99922
rect 85168 94350 85488 94384
rect 85168 94294 85238 94350
rect 85294 94294 85362 94350
rect 85418 94294 85488 94350
rect 85168 94226 85488 94294
rect 85168 94170 85238 94226
rect 85294 94170 85362 94226
rect 85418 94170 85488 94226
rect 85168 94102 85488 94170
rect 85168 94046 85238 94102
rect 85294 94046 85362 94102
rect 85418 94046 85488 94102
rect 85168 93978 85488 94046
rect 85168 93922 85238 93978
rect 85294 93922 85362 93978
rect 85418 93922 85488 93978
rect 85168 93888 85488 93922
rect 93154 94350 93774 111922
rect 93154 94294 93250 94350
rect 93306 94294 93374 94350
rect 93430 94294 93498 94350
rect 93554 94294 93622 94350
rect 93678 94294 93774 94350
rect 93154 94226 93774 94294
rect 93154 94170 93250 94226
rect 93306 94170 93374 94226
rect 93430 94170 93498 94226
rect 93554 94170 93622 94226
rect 93678 94170 93774 94226
rect 93154 94102 93774 94170
rect 93154 94046 93250 94102
rect 93306 94046 93374 94102
rect 93430 94046 93498 94102
rect 93554 94046 93622 94102
rect 93678 94046 93774 94102
rect 93154 93978 93774 94046
rect 93154 93922 93250 93978
rect 93306 93922 93374 93978
rect 93430 93922 93498 93978
rect 93554 93922 93622 93978
rect 93678 93922 93774 93978
rect 78874 82294 78970 82350
rect 79026 82294 79094 82350
rect 79150 82294 79218 82350
rect 79274 82294 79342 82350
rect 79398 82294 79494 82350
rect 78874 82226 79494 82294
rect 78874 82170 78970 82226
rect 79026 82170 79094 82226
rect 79150 82170 79218 82226
rect 79274 82170 79342 82226
rect 79398 82170 79494 82226
rect 78874 82102 79494 82170
rect 78874 82046 78970 82102
rect 79026 82046 79094 82102
rect 79150 82046 79218 82102
rect 79274 82046 79342 82102
rect 79398 82046 79494 82102
rect 78874 81978 79494 82046
rect 78874 81922 78970 81978
rect 79026 81922 79094 81978
rect 79150 81922 79218 81978
rect 79274 81922 79342 81978
rect 79398 81922 79494 81978
rect 78874 64350 79494 81922
rect 85168 76350 85488 76384
rect 85168 76294 85238 76350
rect 85294 76294 85362 76350
rect 85418 76294 85488 76350
rect 85168 76226 85488 76294
rect 85168 76170 85238 76226
rect 85294 76170 85362 76226
rect 85418 76170 85488 76226
rect 85168 76102 85488 76170
rect 85168 76046 85238 76102
rect 85294 76046 85362 76102
rect 85418 76046 85488 76102
rect 85168 75978 85488 76046
rect 85168 75922 85238 75978
rect 85294 75922 85362 75978
rect 85418 75922 85488 75978
rect 85168 75888 85488 75922
rect 93154 76350 93774 93922
rect 93154 76294 93250 76350
rect 93306 76294 93374 76350
rect 93430 76294 93498 76350
rect 93554 76294 93622 76350
rect 93678 76294 93774 76350
rect 93154 76226 93774 76294
rect 93154 76170 93250 76226
rect 93306 76170 93374 76226
rect 93430 76170 93498 76226
rect 93554 76170 93622 76226
rect 93678 76170 93774 76226
rect 93154 76102 93774 76170
rect 93154 76046 93250 76102
rect 93306 76046 93374 76102
rect 93430 76046 93498 76102
rect 93554 76046 93622 76102
rect 93678 76046 93774 76102
rect 93154 75978 93774 76046
rect 93154 75922 93250 75978
rect 93306 75922 93374 75978
rect 93430 75922 93498 75978
rect 93554 75922 93622 75978
rect 93678 75922 93774 75978
rect 78874 64294 78970 64350
rect 79026 64294 79094 64350
rect 79150 64294 79218 64350
rect 79274 64294 79342 64350
rect 79398 64294 79494 64350
rect 78874 64226 79494 64294
rect 78874 64170 78970 64226
rect 79026 64170 79094 64226
rect 79150 64170 79218 64226
rect 79274 64170 79342 64226
rect 79398 64170 79494 64226
rect 78874 64102 79494 64170
rect 78874 64046 78970 64102
rect 79026 64046 79094 64102
rect 79150 64046 79218 64102
rect 79274 64046 79342 64102
rect 79398 64046 79494 64102
rect 78874 63978 79494 64046
rect 78874 63922 78970 63978
rect 79026 63922 79094 63978
rect 79150 63922 79218 63978
rect 79274 63922 79342 63978
rect 79398 63922 79494 63978
rect 78874 46350 79494 63922
rect 85168 58350 85488 58384
rect 85168 58294 85238 58350
rect 85294 58294 85362 58350
rect 85418 58294 85488 58350
rect 85168 58226 85488 58294
rect 85168 58170 85238 58226
rect 85294 58170 85362 58226
rect 85418 58170 85488 58226
rect 85168 58102 85488 58170
rect 85168 58046 85238 58102
rect 85294 58046 85362 58102
rect 85418 58046 85488 58102
rect 85168 57978 85488 58046
rect 85168 57922 85238 57978
rect 85294 57922 85362 57978
rect 85418 57922 85488 57978
rect 85168 57888 85488 57922
rect 93154 58350 93774 75922
rect 93154 58294 93250 58350
rect 93306 58294 93374 58350
rect 93430 58294 93498 58350
rect 93554 58294 93622 58350
rect 93678 58294 93774 58350
rect 93154 58226 93774 58294
rect 93154 58170 93250 58226
rect 93306 58170 93374 58226
rect 93430 58170 93498 58226
rect 93554 58170 93622 58226
rect 93678 58170 93774 58226
rect 93154 58102 93774 58170
rect 93154 58046 93250 58102
rect 93306 58046 93374 58102
rect 93430 58046 93498 58102
rect 93554 58046 93622 58102
rect 93678 58046 93774 58102
rect 93154 57978 93774 58046
rect 93154 57922 93250 57978
rect 93306 57922 93374 57978
rect 93430 57922 93498 57978
rect 93554 57922 93622 57978
rect 93678 57922 93774 57978
rect 78874 46294 78970 46350
rect 79026 46294 79094 46350
rect 79150 46294 79218 46350
rect 79274 46294 79342 46350
rect 79398 46294 79494 46350
rect 78874 46226 79494 46294
rect 78874 46170 78970 46226
rect 79026 46170 79094 46226
rect 79150 46170 79218 46226
rect 79274 46170 79342 46226
rect 79398 46170 79494 46226
rect 78874 46102 79494 46170
rect 78874 46046 78970 46102
rect 79026 46046 79094 46102
rect 79150 46046 79218 46102
rect 79274 46046 79342 46102
rect 79398 46046 79494 46102
rect 78874 45978 79494 46046
rect 78874 45922 78970 45978
rect 79026 45922 79094 45978
rect 79150 45922 79218 45978
rect 79274 45922 79342 45978
rect 79398 45922 79494 45978
rect 78874 28350 79494 45922
rect 85168 40350 85488 40384
rect 85168 40294 85238 40350
rect 85294 40294 85362 40350
rect 85418 40294 85488 40350
rect 85168 40226 85488 40294
rect 85168 40170 85238 40226
rect 85294 40170 85362 40226
rect 85418 40170 85488 40226
rect 85168 40102 85488 40170
rect 85168 40046 85238 40102
rect 85294 40046 85362 40102
rect 85418 40046 85488 40102
rect 85168 39978 85488 40046
rect 85168 39922 85238 39978
rect 85294 39922 85362 39978
rect 85418 39922 85488 39978
rect 85168 39888 85488 39922
rect 93154 40350 93774 57922
rect 93154 40294 93250 40350
rect 93306 40294 93374 40350
rect 93430 40294 93498 40350
rect 93554 40294 93622 40350
rect 93678 40294 93774 40350
rect 93154 40226 93774 40294
rect 93154 40170 93250 40226
rect 93306 40170 93374 40226
rect 93430 40170 93498 40226
rect 93554 40170 93622 40226
rect 93678 40170 93774 40226
rect 93154 40102 93774 40170
rect 93154 40046 93250 40102
rect 93306 40046 93374 40102
rect 93430 40046 93498 40102
rect 93554 40046 93622 40102
rect 93678 40046 93774 40102
rect 93154 39978 93774 40046
rect 93154 39922 93250 39978
rect 93306 39922 93374 39978
rect 93430 39922 93498 39978
rect 93554 39922 93622 39978
rect 93678 39922 93774 39978
rect 78874 28294 78970 28350
rect 79026 28294 79094 28350
rect 79150 28294 79218 28350
rect 79274 28294 79342 28350
rect 79398 28294 79494 28350
rect 78874 28226 79494 28294
rect 78874 28170 78970 28226
rect 79026 28170 79094 28226
rect 79150 28170 79218 28226
rect 79274 28170 79342 28226
rect 79398 28170 79494 28226
rect 78874 28102 79494 28170
rect 78874 28046 78970 28102
rect 79026 28046 79094 28102
rect 79150 28046 79218 28102
rect 79274 28046 79342 28102
rect 79398 28046 79494 28102
rect 78874 27978 79494 28046
rect 78874 27922 78970 27978
rect 79026 27922 79094 27978
rect 79150 27922 79218 27978
rect 79274 27922 79342 27978
rect 79398 27922 79494 27978
rect 78874 10350 79494 27922
rect 78874 10294 78970 10350
rect 79026 10294 79094 10350
rect 79150 10294 79218 10350
rect 79274 10294 79342 10350
rect 79398 10294 79494 10350
rect 78874 10226 79494 10294
rect 78874 10170 78970 10226
rect 79026 10170 79094 10226
rect 79150 10170 79218 10226
rect 79274 10170 79342 10226
rect 79398 10170 79494 10226
rect 78874 10102 79494 10170
rect 78874 10046 78970 10102
rect 79026 10046 79094 10102
rect 79150 10046 79218 10102
rect 79274 10046 79342 10102
rect 79398 10046 79494 10102
rect 78874 9978 79494 10046
rect 78874 9922 78970 9978
rect 79026 9922 79094 9978
rect 79150 9922 79218 9978
rect 79274 9922 79342 9978
rect 79398 9922 79494 9978
rect 78874 -1120 79494 9922
rect 78874 -1176 78970 -1120
rect 79026 -1176 79094 -1120
rect 79150 -1176 79218 -1120
rect 79274 -1176 79342 -1120
rect 79398 -1176 79494 -1120
rect 78874 -1244 79494 -1176
rect 78874 -1300 78970 -1244
rect 79026 -1300 79094 -1244
rect 79150 -1300 79218 -1244
rect 79274 -1300 79342 -1244
rect 79398 -1300 79494 -1244
rect 78874 -1368 79494 -1300
rect 78874 -1424 78970 -1368
rect 79026 -1424 79094 -1368
rect 79150 -1424 79218 -1368
rect 79274 -1424 79342 -1368
rect 79398 -1424 79494 -1368
rect 78874 -1492 79494 -1424
rect 78874 -1548 78970 -1492
rect 79026 -1548 79094 -1492
rect 79150 -1548 79218 -1492
rect 79274 -1548 79342 -1492
rect 79398 -1548 79494 -1492
rect 78874 -1644 79494 -1548
rect 93154 22350 93774 39922
rect 93154 22294 93250 22350
rect 93306 22294 93374 22350
rect 93430 22294 93498 22350
rect 93554 22294 93622 22350
rect 93678 22294 93774 22350
rect 93154 22226 93774 22294
rect 93154 22170 93250 22226
rect 93306 22170 93374 22226
rect 93430 22170 93498 22226
rect 93554 22170 93622 22226
rect 93678 22170 93774 22226
rect 93154 22102 93774 22170
rect 93154 22046 93250 22102
rect 93306 22046 93374 22102
rect 93430 22046 93498 22102
rect 93554 22046 93622 22102
rect 93678 22046 93774 22102
rect 93154 21978 93774 22046
rect 93154 21922 93250 21978
rect 93306 21922 93374 21978
rect 93430 21922 93498 21978
rect 93554 21922 93622 21978
rect 93678 21922 93774 21978
rect 93154 4350 93774 21922
rect 93154 4294 93250 4350
rect 93306 4294 93374 4350
rect 93430 4294 93498 4350
rect 93554 4294 93622 4350
rect 93678 4294 93774 4350
rect 93154 4226 93774 4294
rect 93154 4170 93250 4226
rect 93306 4170 93374 4226
rect 93430 4170 93498 4226
rect 93554 4170 93622 4226
rect 93678 4170 93774 4226
rect 93154 4102 93774 4170
rect 93154 4046 93250 4102
rect 93306 4046 93374 4102
rect 93430 4046 93498 4102
rect 93554 4046 93622 4102
rect 93678 4046 93774 4102
rect 93154 3978 93774 4046
rect 93154 3922 93250 3978
rect 93306 3922 93374 3978
rect 93430 3922 93498 3978
rect 93554 3922 93622 3978
rect 93678 3922 93774 3978
rect 93154 -160 93774 3922
rect 93154 -216 93250 -160
rect 93306 -216 93374 -160
rect 93430 -216 93498 -160
rect 93554 -216 93622 -160
rect 93678 -216 93774 -160
rect 93154 -284 93774 -216
rect 93154 -340 93250 -284
rect 93306 -340 93374 -284
rect 93430 -340 93498 -284
rect 93554 -340 93622 -284
rect 93678 -340 93774 -284
rect 93154 -408 93774 -340
rect 93154 -464 93250 -408
rect 93306 -464 93374 -408
rect 93430 -464 93498 -408
rect 93554 -464 93622 -408
rect 93678 -464 93774 -408
rect 93154 -532 93774 -464
rect 93154 -588 93250 -532
rect 93306 -588 93374 -532
rect 93430 -588 93498 -532
rect 93554 -588 93622 -532
rect 93678 -588 93774 -532
rect 93154 -1644 93774 -588
rect 96874 598172 97494 598268
rect 96874 598116 96970 598172
rect 97026 598116 97094 598172
rect 97150 598116 97218 598172
rect 97274 598116 97342 598172
rect 97398 598116 97494 598172
rect 96874 598048 97494 598116
rect 96874 597992 96970 598048
rect 97026 597992 97094 598048
rect 97150 597992 97218 598048
rect 97274 597992 97342 598048
rect 97398 597992 97494 598048
rect 96874 597924 97494 597992
rect 96874 597868 96970 597924
rect 97026 597868 97094 597924
rect 97150 597868 97218 597924
rect 97274 597868 97342 597924
rect 97398 597868 97494 597924
rect 96874 597800 97494 597868
rect 96874 597744 96970 597800
rect 97026 597744 97094 597800
rect 97150 597744 97218 597800
rect 97274 597744 97342 597800
rect 97398 597744 97494 597800
rect 96874 586350 97494 597744
rect 96874 586294 96970 586350
rect 97026 586294 97094 586350
rect 97150 586294 97218 586350
rect 97274 586294 97342 586350
rect 97398 586294 97494 586350
rect 96874 586226 97494 586294
rect 96874 586170 96970 586226
rect 97026 586170 97094 586226
rect 97150 586170 97218 586226
rect 97274 586170 97342 586226
rect 97398 586170 97494 586226
rect 96874 586102 97494 586170
rect 96874 586046 96970 586102
rect 97026 586046 97094 586102
rect 97150 586046 97218 586102
rect 97274 586046 97342 586102
rect 97398 586046 97494 586102
rect 96874 585978 97494 586046
rect 96874 585922 96970 585978
rect 97026 585922 97094 585978
rect 97150 585922 97218 585978
rect 97274 585922 97342 585978
rect 97398 585922 97494 585978
rect 96874 568350 97494 585922
rect 96874 568294 96970 568350
rect 97026 568294 97094 568350
rect 97150 568294 97218 568350
rect 97274 568294 97342 568350
rect 97398 568294 97494 568350
rect 96874 568226 97494 568294
rect 96874 568170 96970 568226
rect 97026 568170 97094 568226
rect 97150 568170 97218 568226
rect 97274 568170 97342 568226
rect 97398 568170 97494 568226
rect 96874 568102 97494 568170
rect 96874 568046 96970 568102
rect 97026 568046 97094 568102
rect 97150 568046 97218 568102
rect 97274 568046 97342 568102
rect 97398 568046 97494 568102
rect 96874 567978 97494 568046
rect 96874 567922 96970 567978
rect 97026 567922 97094 567978
rect 97150 567922 97218 567978
rect 97274 567922 97342 567978
rect 97398 567922 97494 567978
rect 96874 550350 97494 567922
rect 96874 550294 96970 550350
rect 97026 550294 97094 550350
rect 97150 550294 97218 550350
rect 97274 550294 97342 550350
rect 97398 550294 97494 550350
rect 96874 550226 97494 550294
rect 96874 550170 96970 550226
rect 97026 550170 97094 550226
rect 97150 550170 97218 550226
rect 97274 550170 97342 550226
rect 97398 550170 97494 550226
rect 96874 550102 97494 550170
rect 96874 550046 96970 550102
rect 97026 550046 97094 550102
rect 97150 550046 97218 550102
rect 97274 550046 97342 550102
rect 97398 550046 97494 550102
rect 96874 549978 97494 550046
rect 96874 549922 96970 549978
rect 97026 549922 97094 549978
rect 97150 549922 97218 549978
rect 97274 549922 97342 549978
rect 97398 549922 97494 549978
rect 96874 532350 97494 549922
rect 96874 532294 96970 532350
rect 97026 532294 97094 532350
rect 97150 532294 97218 532350
rect 97274 532294 97342 532350
rect 97398 532294 97494 532350
rect 96874 532226 97494 532294
rect 96874 532170 96970 532226
rect 97026 532170 97094 532226
rect 97150 532170 97218 532226
rect 97274 532170 97342 532226
rect 97398 532170 97494 532226
rect 96874 532102 97494 532170
rect 96874 532046 96970 532102
rect 97026 532046 97094 532102
rect 97150 532046 97218 532102
rect 97274 532046 97342 532102
rect 97398 532046 97494 532102
rect 96874 531978 97494 532046
rect 96874 531922 96970 531978
rect 97026 531922 97094 531978
rect 97150 531922 97218 531978
rect 97274 531922 97342 531978
rect 97398 531922 97494 531978
rect 96874 514350 97494 531922
rect 111154 597212 111774 598268
rect 111154 597156 111250 597212
rect 111306 597156 111374 597212
rect 111430 597156 111498 597212
rect 111554 597156 111622 597212
rect 111678 597156 111774 597212
rect 111154 597088 111774 597156
rect 111154 597032 111250 597088
rect 111306 597032 111374 597088
rect 111430 597032 111498 597088
rect 111554 597032 111622 597088
rect 111678 597032 111774 597088
rect 111154 596964 111774 597032
rect 111154 596908 111250 596964
rect 111306 596908 111374 596964
rect 111430 596908 111498 596964
rect 111554 596908 111622 596964
rect 111678 596908 111774 596964
rect 111154 596840 111774 596908
rect 111154 596784 111250 596840
rect 111306 596784 111374 596840
rect 111430 596784 111498 596840
rect 111554 596784 111622 596840
rect 111678 596784 111774 596840
rect 111154 580350 111774 596784
rect 111154 580294 111250 580350
rect 111306 580294 111374 580350
rect 111430 580294 111498 580350
rect 111554 580294 111622 580350
rect 111678 580294 111774 580350
rect 111154 580226 111774 580294
rect 111154 580170 111250 580226
rect 111306 580170 111374 580226
rect 111430 580170 111498 580226
rect 111554 580170 111622 580226
rect 111678 580170 111774 580226
rect 111154 580102 111774 580170
rect 111154 580046 111250 580102
rect 111306 580046 111374 580102
rect 111430 580046 111498 580102
rect 111554 580046 111622 580102
rect 111678 580046 111774 580102
rect 111154 579978 111774 580046
rect 111154 579922 111250 579978
rect 111306 579922 111374 579978
rect 111430 579922 111498 579978
rect 111554 579922 111622 579978
rect 111678 579922 111774 579978
rect 111154 562350 111774 579922
rect 111154 562294 111250 562350
rect 111306 562294 111374 562350
rect 111430 562294 111498 562350
rect 111554 562294 111622 562350
rect 111678 562294 111774 562350
rect 111154 562226 111774 562294
rect 111154 562170 111250 562226
rect 111306 562170 111374 562226
rect 111430 562170 111498 562226
rect 111554 562170 111622 562226
rect 111678 562170 111774 562226
rect 111154 562102 111774 562170
rect 111154 562046 111250 562102
rect 111306 562046 111374 562102
rect 111430 562046 111498 562102
rect 111554 562046 111622 562102
rect 111678 562046 111774 562102
rect 111154 561978 111774 562046
rect 111154 561922 111250 561978
rect 111306 561922 111374 561978
rect 111430 561922 111498 561978
rect 111554 561922 111622 561978
rect 111678 561922 111774 561978
rect 111154 544350 111774 561922
rect 111154 544294 111250 544350
rect 111306 544294 111374 544350
rect 111430 544294 111498 544350
rect 111554 544294 111622 544350
rect 111678 544294 111774 544350
rect 111154 544226 111774 544294
rect 111154 544170 111250 544226
rect 111306 544170 111374 544226
rect 111430 544170 111498 544226
rect 111554 544170 111622 544226
rect 111678 544170 111774 544226
rect 111154 544102 111774 544170
rect 111154 544046 111250 544102
rect 111306 544046 111374 544102
rect 111430 544046 111498 544102
rect 111554 544046 111622 544102
rect 111678 544046 111774 544102
rect 111154 543978 111774 544046
rect 111154 543922 111250 543978
rect 111306 543922 111374 543978
rect 111430 543922 111498 543978
rect 111554 543922 111622 543978
rect 111678 543922 111774 543978
rect 111154 526350 111774 543922
rect 114874 598172 115494 598268
rect 114874 598116 114970 598172
rect 115026 598116 115094 598172
rect 115150 598116 115218 598172
rect 115274 598116 115342 598172
rect 115398 598116 115494 598172
rect 114874 598048 115494 598116
rect 114874 597992 114970 598048
rect 115026 597992 115094 598048
rect 115150 597992 115218 598048
rect 115274 597992 115342 598048
rect 115398 597992 115494 598048
rect 114874 597924 115494 597992
rect 114874 597868 114970 597924
rect 115026 597868 115094 597924
rect 115150 597868 115218 597924
rect 115274 597868 115342 597924
rect 115398 597868 115494 597924
rect 114874 597800 115494 597868
rect 114874 597744 114970 597800
rect 115026 597744 115094 597800
rect 115150 597744 115218 597800
rect 115274 597744 115342 597800
rect 115398 597744 115494 597800
rect 114874 586350 115494 597744
rect 114874 586294 114970 586350
rect 115026 586294 115094 586350
rect 115150 586294 115218 586350
rect 115274 586294 115342 586350
rect 115398 586294 115494 586350
rect 114874 586226 115494 586294
rect 114874 586170 114970 586226
rect 115026 586170 115094 586226
rect 115150 586170 115218 586226
rect 115274 586170 115342 586226
rect 115398 586170 115494 586226
rect 114874 586102 115494 586170
rect 114874 586046 114970 586102
rect 115026 586046 115094 586102
rect 115150 586046 115218 586102
rect 115274 586046 115342 586102
rect 115398 586046 115494 586102
rect 114874 585978 115494 586046
rect 114874 585922 114970 585978
rect 115026 585922 115094 585978
rect 115150 585922 115218 585978
rect 115274 585922 115342 585978
rect 115398 585922 115494 585978
rect 114874 568350 115494 585922
rect 114874 568294 114970 568350
rect 115026 568294 115094 568350
rect 115150 568294 115218 568350
rect 115274 568294 115342 568350
rect 115398 568294 115494 568350
rect 114874 568226 115494 568294
rect 114874 568170 114970 568226
rect 115026 568170 115094 568226
rect 115150 568170 115218 568226
rect 115274 568170 115342 568226
rect 115398 568170 115494 568226
rect 114874 568102 115494 568170
rect 114874 568046 114970 568102
rect 115026 568046 115094 568102
rect 115150 568046 115218 568102
rect 115274 568046 115342 568102
rect 115398 568046 115494 568102
rect 114874 567978 115494 568046
rect 114874 567922 114970 567978
rect 115026 567922 115094 567978
rect 115150 567922 115218 567978
rect 115274 567922 115342 567978
rect 115398 567922 115494 567978
rect 114874 550350 115494 567922
rect 114874 550294 114970 550350
rect 115026 550294 115094 550350
rect 115150 550294 115218 550350
rect 115274 550294 115342 550350
rect 115398 550294 115494 550350
rect 114874 550226 115494 550294
rect 114874 550170 114970 550226
rect 115026 550170 115094 550226
rect 115150 550170 115218 550226
rect 115274 550170 115342 550226
rect 115398 550170 115494 550226
rect 114874 550102 115494 550170
rect 114874 550046 114970 550102
rect 115026 550046 115094 550102
rect 115150 550046 115218 550102
rect 115274 550046 115342 550102
rect 115398 550046 115494 550102
rect 114874 549978 115494 550046
rect 114874 549922 114970 549978
rect 115026 549922 115094 549978
rect 115150 549922 115218 549978
rect 115274 549922 115342 549978
rect 115398 549922 115494 549978
rect 114874 532350 115494 549922
rect 114874 532294 114970 532350
rect 115026 532294 115094 532350
rect 115150 532294 115218 532350
rect 115274 532294 115342 532350
rect 115398 532294 115494 532350
rect 114874 532226 115494 532294
rect 114874 532170 114970 532226
rect 115026 532170 115094 532226
rect 115150 532170 115218 532226
rect 115274 532170 115342 532226
rect 115398 532170 115494 532226
rect 114874 532102 115494 532170
rect 114874 532046 114970 532102
rect 115026 532046 115094 532102
rect 115150 532046 115218 532102
rect 115274 532046 115342 532102
rect 115398 532046 115494 532102
rect 114874 531978 115494 532046
rect 114874 531922 114970 531978
rect 115026 531922 115094 531978
rect 115150 531922 115218 531978
rect 115274 531922 115342 531978
rect 115398 531922 115494 531978
rect 114874 527750 115494 531922
rect 129154 597212 129774 598268
rect 129154 597156 129250 597212
rect 129306 597156 129374 597212
rect 129430 597156 129498 597212
rect 129554 597156 129622 597212
rect 129678 597156 129774 597212
rect 129154 597088 129774 597156
rect 129154 597032 129250 597088
rect 129306 597032 129374 597088
rect 129430 597032 129498 597088
rect 129554 597032 129622 597088
rect 129678 597032 129774 597088
rect 129154 596964 129774 597032
rect 129154 596908 129250 596964
rect 129306 596908 129374 596964
rect 129430 596908 129498 596964
rect 129554 596908 129622 596964
rect 129678 596908 129774 596964
rect 129154 596840 129774 596908
rect 129154 596784 129250 596840
rect 129306 596784 129374 596840
rect 129430 596784 129498 596840
rect 129554 596784 129622 596840
rect 129678 596784 129774 596840
rect 129154 580350 129774 596784
rect 129154 580294 129250 580350
rect 129306 580294 129374 580350
rect 129430 580294 129498 580350
rect 129554 580294 129622 580350
rect 129678 580294 129774 580350
rect 129154 580226 129774 580294
rect 129154 580170 129250 580226
rect 129306 580170 129374 580226
rect 129430 580170 129498 580226
rect 129554 580170 129622 580226
rect 129678 580170 129774 580226
rect 129154 580102 129774 580170
rect 129154 580046 129250 580102
rect 129306 580046 129374 580102
rect 129430 580046 129498 580102
rect 129554 580046 129622 580102
rect 129678 580046 129774 580102
rect 129154 579978 129774 580046
rect 129154 579922 129250 579978
rect 129306 579922 129374 579978
rect 129430 579922 129498 579978
rect 129554 579922 129622 579978
rect 129678 579922 129774 579978
rect 129154 562350 129774 579922
rect 129154 562294 129250 562350
rect 129306 562294 129374 562350
rect 129430 562294 129498 562350
rect 129554 562294 129622 562350
rect 129678 562294 129774 562350
rect 129154 562226 129774 562294
rect 129154 562170 129250 562226
rect 129306 562170 129374 562226
rect 129430 562170 129498 562226
rect 129554 562170 129622 562226
rect 129678 562170 129774 562226
rect 129154 562102 129774 562170
rect 129154 562046 129250 562102
rect 129306 562046 129374 562102
rect 129430 562046 129498 562102
rect 129554 562046 129622 562102
rect 129678 562046 129774 562102
rect 129154 561978 129774 562046
rect 129154 561922 129250 561978
rect 129306 561922 129374 561978
rect 129430 561922 129498 561978
rect 129554 561922 129622 561978
rect 129678 561922 129774 561978
rect 129154 544350 129774 561922
rect 129154 544294 129250 544350
rect 129306 544294 129374 544350
rect 129430 544294 129498 544350
rect 129554 544294 129622 544350
rect 129678 544294 129774 544350
rect 129154 544226 129774 544294
rect 129154 544170 129250 544226
rect 129306 544170 129374 544226
rect 129430 544170 129498 544226
rect 129554 544170 129622 544226
rect 129678 544170 129774 544226
rect 129154 544102 129774 544170
rect 129154 544046 129250 544102
rect 129306 544046 129374 544102
rect 129430 544046 129498 544102
rect 129554 544046 129622 544102
rect 129678 544046 129774 544102
rect 129154 543978 129774 544046
rect 129154 543922 129250 543978
rect 129306 543922 129374 543978
rect 129430 543922 129498 543978
rect 129554 543922 129622 543978
rect 129678 543922 129774 543978
rect 129154 527750 129774 543922
rect 132874 598172 133494 598268
rect 132874 598116 132970 598172
rect 133026 598116 133094 598172
rect 133150 598116 133218 598172
rect 133274 598116 133342 598172
rect 133398 598116 133494 598172
rect 132874 598048 133494 598116
rect 132874 597992 132970 598048
rect 133026 597992 133094 598048
rect 133150 597992 133218 598048
rect 133274 597992 133342 598048
rect 133398 597992 133494 598048
rect 132874 597924 133494 597992
rect 132874 597868 132970 597924
rect 133026 597868 133094 597924
rect 133150 597868 133218 597924
rect 133274 597868 133342 597924
rect 133398 597868 133494 597924
rect 132874 597800 133494 597868
rect 132874 597744 132970 597800
rect 133026 597744 133094 597800
rect 133150 597744 133218 597800
rect 133274 597744 133342 597800
rect 133398 597744 133494 597800
rect 132874 586350 133494 597744
rect 132874 586294 132970 586350
rect 133026 586294 133094 586350
rect 133150 586294 133218 586350
rect 133274 586294 133342 586350
rect 133398 586294 133494 586350
rect 132874 586226 133494 586294
rect 132874 586170 132970 586226
rect 133026 586170 133094 586226
rect 133150 586170 133218 586226
rect 133274 586170 133342 586226
rect 133398 586170 133494 586226
rect 132874 586102 133494 586170
rect 132874 586046 132970 586102
rect 133026 586046 133094 586102
rect 133150 586046 133218 586102
rect 133274 586046 133342 586102
rect 133398 586046 133494 586102
rect 132874 585978 133494 586046
rect 132874 585922 132970 585978
rect 133026 585922 133094 585978
rect 133150 585922 133218 585978
rect 133274 585922 133342 585978
rect 133398 585922 133494 585978
rect 132874 568350 133494 585922
rect 132874 568294 132970 568350
rect 133026 568294 133094 568350
rect 133150 568294 133218 568350
rect 133274 568294 133342 568350
rect 133398 568294 133494 568350
rect 132874 568226 133494 568294
rect 132874 568170 132970 568226
rect 133026 568170 133094 568226
rect 133150 568170 133218 568226
rect 133274 568170 133342 568226
rect 133398 568170 133494 568226
rect 132874 568102 133494 568170
rect 132874 568046 132970 568102
rect 133026 568046 133094 568102
rect 133150 568046 133218 568102
rect 133274 568046 133342 568102
rect 133398 568046 133494 568102
rect 132874 567978 133494 568046
rect 132874 567922 132970 567978
rect 133026 567922 133094 567978
rect 133150 567922 133218 567978
rect 133274 567922 133342 567978
rect 133398 567922 133494 567978
rect 132874 550350 133494 567922
rect 132874 550294 132970 550350
rect 133026 550294 133094 550350
rect 133150 550294 133218 550350
rect 133274 550294 133342 550350
rect 133398 550294 133494 550350
rect 132874 550226 133494 550294
rect 132874 550170 132970 550226
rect 133026 550170 133094 550226
rect 133150 550170 133218 550226
rect 133274 550170 133342 550226
rect 133398 550170 133494 550226
rect 132874 550102 133494 550170
rect 132874 550046 132970 550102
rect 133026 550046 133094 550102
rect 133150 550046 133218 550102
rect 133274 550046 133342 550102
rect 133398 550046 133494 550102
rect 132874 549978 133494 550046
rect 132874 549922 132970 549978
rect 133026 549922 133094 549978
rect 133150 549922 133218 549978
rect 133274 549922 133342 549978
rect 133398 549922 133494 549978
rect 132874 532350 133494 549922
rect 132874 532294 132970 532350
rect 133026 532294 133094 532350
rect 133150 532294 133218 532350
rect 133274 532294 133342 532350
rect 133398 532294 133494 532350
rect 132874 532226 133494 532294
rect 132874 532170 132970 532226
rect 133026 532170 133094 532226
rect 133150 532170 133218 532226
rect 133274 532170 133342 532226
rect 133398 532170 133494 532226
rect 132874 532102 133494 532170
rect 132874 532046 132970 532102
rect 133026 532046 133094 532102
rect 133150 532046 133218 532102
rect 133274 532046 133342 532102
rect 133398 532046 133494 532102
rect 132874 531978 133494 532046
rect 132874 531922 132970 531978
rect 133026 531922 133094 531978
rect 133150 531922 133218 531978
rect 133274 531922 133342 531978
rect 133398 531922 133494 531978
rect 132874 527750 133494 531922
rect 147154 597212 147774 598268
rect 147154 597156 147250 597212
rect 147306 597156 147374 597212
rect 147430 597156 147498 597212
rect 147554 597156 147622 597212
rect 147678 597156 147774 597212
rect 147154 597088 147774 597156
rect 147154 597032 147250 597088
rect 147306 597032 147374 597088
rect 147430 597032 147498 597088
rect 147554 597032 147622 597088
rect 147678 597032 147774 597088
rect 147154 596964 147774 597032
rect 147154 596908 147250 596964
rect 147306 596908 147374 596964
rect 147430 596908 147498 596964
rect 147554 596908 147622 596964
rect 147678 596908 147774 596964
rect 147154 596840 147774 596908
rect 147154 596784 147250 596840
rect 147306 596784 147374 596840
rect 147430 596784 147498 596840
rect 147554 596784 147622 596840
rect 147678 596784 147774 596840
rect 147154 580350 147774 596784
rect 147154 580294 147250 580350
rect 147306 580294 147374 580350
rect 147430 580294 147498 580350
rect 147554 580294 147622 580350
rect 147678 580294 147774 580350
rect 147154 580226 147774 580294
rect 147154 580170 147250 580226
rect 147306 580170 147374 580226
rect 147430 580170 147498 580226
rect 147554 580170 147622 580226
rect 147678 580170 147774 580226
rect 147154 580102 147774 580170
rect 147154 580046 147250 580102
rect 147306 580046 147374 580102
rect 147430 580046 147498 580102
rect 147554 580046 147622 580102
rect 147678 580046 147774 580102
rect 147154 579978 147774 580046
rect 147154 579922 147250 579978
rect 147306 579922 147374 579978
rect 147430 579922 147498 579978
rect 147554 579922 147622 579978
rect 147678 579922 147774 579978
rect 147154 562350 147774 579922
rect 147154 562294 147250 562350
rect 147306 562294 147374 562350
rect 147430 562294 147498 562350
rect 147554 562294 147622 562350
rect 147678 562294 147774 562350
rect 147154 562226 147774 562294
rect 147154 562170 147250 562226
rect 147306 562170 147374 562226
rect 147430 562170 147498 562226
rect 147554 562170 147622 562226
rect 147678 562170 147774 562226
rect 147154 562102 147774 562170
rect 147154 562046 147250 562102
rect 147306 562046 147374 562102
rect 147430 562046 147498 562102
rect 147554 562046 147622 562102
rect 147678 562046 147774 562102
rect 147154 561978 147774 562046
rect 147154 561922 147250 561978
rect 147306 561922 147374 561978
rect 147430 561922 147498 561978
rect 147554 561922 147622 561978
rect 147678 561922 147774 561978
rect 147154 544350 147774 561922
rect 147154 544294 147250 544350
rect 147306 544294 147374 544350
rect 147430 544294 147498 544350
rect 147554 544294 147622 544350
rect 147678 544294 147774 544350
rect 147154 544226 147774 544294
rect 147154 544170 147250 544226
rect 147306 544170 147374 544226
rect 147430 544170 147498 544226
rect 147554 544170 147622 544226
rect 147678 544170 147774 544226
rect 147154 544102 147774 544170
rect 147154 544046 147250 544102
rect 147306 544046 147374 544102
rect 147430 544046 147498 544102
rect 147554 544046 147622 544102
rect 147678 544046 147774 544102
rect 147154 543978 147774 544046
rect 147154 543922 147250 543978
rect 147306 543922 147374 543978
rect 147430 543922 147498 543978
rect 147554 543922 147622 543978
rect 147678 543922 147774 543978
rect 147154 527750 147774 543922
rect 150874 598172 151494 598268
rect 150874 598116 150970 598172
rect 151026 598116 151094 598172
rect 151150 598116 151218 598172
rect 151274 598116 151342 598172
rect 151398 598116 151494 598172
rect 150874 598048 151494 598116
rect 150874 597992 150970 598048
rect 151026 597992 151094 598048
rect 151150 597992 151218 598048
rect 151274 597992 151342 598048
rect 151398 597992 151494 598048
rect 150874 597924 151494 597992
rect 150874 597868 150970 597924
rect 151026 597868 151094 597924
rect 151150 597868 151218 597924
rect 151274 597868 151342 597924
rect 151398 597868 151494 597924
rect 150874 597800 151494 597868
rect 150874 597744 150970 597800
rect 151026 597744 151094 597800
rect 151150 597744 151218 597800
rect 151274 597744 151342 597800
rect 151398 597744 151494 597800
rect 150874 586350 151494 597744
rect 150874 586294 150970 586350
rect 151026 586294 151094 586350
rect 151150 586294 151218 586350
rect 151274 586294 151342 586350
rect 151398 586294 151494 586350
rect 150874 586226 151494 586294
rect 150874 586170 150970 586226
rect 151026 586170 151094 586226
rect 151150 586170 151218 586226
rect 151274 586170 151342 586226
rect 151398 586170 151494 586226
rect 150874 586102 151494 586170
rect 150874 586046 150970 586102
rect 151026 586046 151094 586102
rect 151150 586046 151218 586102
rect 151274 586046 151342 586102
rect 151398 586046 151494 586102
rect 150874 585978 151494 586046
rect 150874 585922 150970 585978
rect 151026 585922 151094 585978
rect 151150 585922 151218 585978
rect 151274 585922 151342 585978
rect 151398 585922 151494 585978
rect 150874 568350 151494 585922
rect 150874 568294 150970 568350
rect 151026 568294 151094 568350
rect 151150 568294 151218 568350
rect 151274 568294 151342 568350
rect 151398 568294 151494 568350
rect 150874 568226 151494 568294
rect 150874 568170 150970 568226
rect 151026 568170 151094 568226
rect 151150 568170 151218 568226
rect 151274 568170 151342 568226
rect 151398 568170 151494 568226
rect 150874 568102 151494 568170
rect 150874 568046 150970 568102
rect 151026 568046 151094 568102
rect 151150 568046 151218 568102
rect 151274 568046 151342 568102
rect 151398 568046 151494 568102
rect 150874 567978 151494 568046
rect 150874 567922 150970 567978
rect 151026 567922 151094 567978
rect 151150 567922 151218 567978
rect 151274 567922 151342 567978
rect 151398 567922 151494 567978
rect 150874 550350 151494 567922
rect 150874 550294 150970 550350
rect 151026 550294 151094 550350
rect 151150 550294 151218 550350
rect 151274 550294 151342 550350
rect 151398 550294 151494 550350
rect 150874 550226 151494 550294
rect 150874 550170 150970 550226
rect 151026 550170 151094 550226
rect 151150 550170 151218 550226
rect 151274 550170 151342 550226
rect 151398 550170 151494 550226
rect 150874 550102 151494 550170
rect 150874 550046 150970 550102
rect 151026 550046 151094 550102
rect 151150 550046 151218 550102
rect 151274 550046 151342 550102
rect 151398 550046 151494 550102
rect 150874 549978 151494 550046
rect 150874 549922 150970 549978
rect 151026 549922 151094 549978
rect 151150 549922 151218 549978
rect 151274 549922 151342 549978
rect 151398 549922 151494 549978
rect 150874 532350 151494 549922
rect 150874 532294 150970 532350
rect 151026 532294 151094 532350
rect 151150 532294 151218 532350
rect 151274 532294 151342 532350
rect 151398 532294 151494 532350
rect 150874 532226 151494 532294
rect 150874 532170 150970 532226
rect 151026 532170 151094 532226
rect 151150 532170 151218 532226
rect 151274 532170 151342 532226
rect 151398 532170 151494 532226
rect 150874 532102 151494 532170
rect 150874 532046 150970 532102
rect 151026 532046 151094 532102
rect 151150 532046 151218 532102
rect 151274 532046 151342 532102
rect 151398 532046 151494 532102
rect 150874 531978 151494 532046
rect 150874 531922 150970 531978
rect 151026 531922 151094 531978
rect 151150 531922 151218 531978
rect 151274 531922 151342 531978
rect 151398 531922 151494 531978
rect 150874 527750 151494 531922
rect 165154 597212 165774 598268
rect 165154 597156 165250 597212
rect 165306 597156 165374 597212
rect 165430 597156 165498 597212
rect 165554 597156 165622 597212
rect 165678 597156 165774 597212
rect 165154 597088 165774 597156
rect 165154 597032 165250 597088
rect 165306 597032 165374 597088
rect 165430 597032 165498 597088
rect 165554 597032 165622 597088
rect 165678 597032 165774 597088
rect 165154 596964 165774 597032
rect 165154 596908 165250 596964
rect 165306 596908 165374 596964
rect 165430 596908 165498 596964
rect 165554 596908 165622 596964
rect 165678 596908 165774 596964
rect 165154 596840 165774 596908
rect 165154 596784 165250 596840
rect 165306 596784 165374 596840
rect 165430 596784 165498 596840
rect 165554 596784 165622 596840
rect 165678 596784 165774 596840
rect 165154 580350 165774 596784
rect 165154 580294 165250 580350
rect 165306 580294 165374 580350
rect 165430 580294 165498 580350
rect 165554 580294 165622 580350
rect 165678 580294 165774 580350
rect 165154 580226 165774 580294
rect 165154 580170 165250 580226
rect 165306 580170 165374 580226
rect 165430 580170 165498 580226
rect 165554 580170 165622 580226
rect 165678 580170 165774 580226
rect 165154 580102 165774 580170
rect 165154 580046 165250 580102
rect 165306 580046 165374 580102
rect 165430 580046 165498 580102
rect 165554 580046 165622 580102
rect 165678 580046 165774 580102
rect 165154 579978 165774 580046
rect 165154 579922 165250 579978
rect 165306 579922 165374 579978
rect 165430 579922 165498 579978
rect 165554 579922 165622 579978
rect 165678 579922 165774 579978
rect 165154 562350 165774 579922
rect 165154 562294 165250 562350
rect 165306 562294 165374 562350
rect 165430 562294 165498 562350
rect 165554 562294 165622 562350
rect 165678 562294 165774 562350
rect 165154 562226 165774 562294
rect 165154 562170 165250 562226
rect 165306 562170 165374 562226
rect 165430 562170 165498 562226
rect 165554 562170 165622 562226
rect 165678 562170 165774 562226
rect 165154 562102 165774 562170
rect 165154 562046 165250 562102
rect 165306 562046 165374 562102
rect 165430 562046 165498 562102
rect 165554 562046 165622 562102
rect 165678 562046 165774 562102
rect 165154 561978 165774 562046
rect 165154 561922 165250 561978
rect 165306 561922 165374 561978
rect 165430 561922 165498 561978
rect 165554 561922 165622 561978
rect 165678 561922 165774 561978
rect 165154 544350 165774 561922
rect 165154 544294 165250 544350
rect 165306 544294 165374 544350
rect 165430 544294 165498 544350
rect 165554 544294 165622 544350
rect 165678 544294 165774 544350
rect 165154 544226 165774 544294
rect 165154 544170 165250 544226
rect 165306 544170 165374 544226
rect 165430 544170 165498 544226
rect 165554 544170 165622 544226
rect 165678 544170 165774 544226
rect 165154 544102 165774 544170
rect 165154 544046 165250 544102
rect 165306 544046 165374 544102
rect 165430 544046 165498 544102
rect 165554 544046 165622 544102
rect 165678 544046 165774 544102
rect 165154 543978 165774 544046
rect 165154 543922 165250 543978
rect 165306 543922 165374 543978
rect 165430 543922 165498 543978
rect 165554 543922 165622 543978
rect 165678 543922 165774 543978
rect 165154 527750 165774 543922
rect 168874 598172 169494 598268
rect 168874 598116 168970 598172
rect 169026 598116 169094 598172
rect 169150 598116 169218 598172
rect 169274 598116 169342 598172
rect 169398 598116 169494 598172
rect 168874 598048 169494 598116
rect 168874 597992 168970 598048
rect 169026 597992 169094 598048
rect 169150 597992 169218 598048
rect 169274 597992 169342 598048
rect 169398 597992 169494 598048
rect 168874 597924 169494 597992
rect 168874 597868 168970 597924
rect 169026 597868 169094 597924
rect 169150 597868 169218 597924
rect 169274 597868 169342 597924
rect 169398 597868 169494 597924
rect 168874 597800 169494 597868
rect 168874 597744 168970 597800
rect 169026 597744 169094 597800
rect 169150 597744 169218 597800
rect 169274 597744 169342 597800
rect 169398 597744 169494 597800
rect 168874 586350 169494 597744
rect 168874 586294 168970 586350
rect 169026 586294 169094 586350
rect 169150 586294 169218 586350
rect 169274 586294 169342 586350
rect 169398 586294 169494 586350
rect 168874 586226 169494 586294
rect 168874 586170 168970 586226
rect 169026 586170 169094 586226
rect 169150 586170 169218 586226
rect 169274 586170 169342 586226
rect 169398 586170 169494 586226
rect 168874 586102 169494 586170
rect 168874 586046 168970 586102
rect 169026 586046 169094 586102
rect 169150 586046 169218 586102
rect 169274 586046 169342 586102
rect 169398 586046 169494 586102
rect 168874 585978 169494 586046
rect 168874 585922 168970 585978
rect 169026 585922 169094 585978
rect 169150 585922 169218 585978
rect 169274 585922 169342 585978
rect 169398 585922 169494 585978
rect 168874 568350 169494 585922
rect 168874 568294 168970 568350
rect 169026 568294 169094 568350
rect 169150 568294 169218 568350
rect 169274 568294 169342 568350
rect 169398 568294 169494 568350
rect 168874 568226 169494 568294
rect 168874 568170 168970 568226
rect 169026 568170 169094 568226
rect 169150 568170 169218 568226
rect 169274 568170 169342 568226
rect 169398 568170 169494 568226
rect 168874 568102 169494 568170
rect 168874 568046 168970 568102
rect 169026 568046 169094 568102
rect 169150 568046 169218 568102
rect 169274 568046 169342 568102
rect 169398 568046 169494 568102
rect 168874 567978 169494 568046
rect 168874 567922 168970 567978
rect 169026 567922 169094 567978
rect 169150 567922 169218 567978
rect 169274 567922 169342 567978
rect 169398 567922 169494 567978
rect 168874 550350 169494 567922
rect 168874 550294 168970 550350
rect 169026 550294 169094 550350
rect 169150 550294 169218 550350
rect 169274 550294 169342 550350
rect 169398 550294 169494 550350
rect 168874 550226 169494 550294
rect 168874 550170 168970 550226
rect 169026 550170 169094 550226
rect 169150 550170 169218 550226
rect 169274 550170 169342 550226
rect 169398 550170 169494 550226
rect 168874 550102 169494 550170
rect 168874 550046 168970 550102
rect 169026 550046 169094 550102
rect 169150 550046 169218 550102
rect 169274 550046 169342 550102
rect 169398 550046 169494 550102
rect 168874 549978 169494 550046
rect 168874 549922 168970 549978
rect 169026 549922 169094 549978
rect 169150 549922 169218 549978
rect 169274 549922 169342 549978
rect 169398 549922 169494 549978
rect 168874 532350 169494 549922
rect 168874 532294 168970 532350
rect 169026 532294 169094 532350
rect 169150 532294 169218 532350
rect 169274 532294 169342 532350
rect 169398 532294 169494 532350
rect 168874 532226 169494 532294
rect 168874 532170 168970 532226
rect 169026 532170 169094 532226
rect 169150 532170 169218 532226
rect 169274 532170 169342 532226
rect 169398 532170 169494 532226
rect 168874 532102 169494 532170
rect 168874 532046 168970 532102
rect 169026 532046 169094 532102
rect 169150 532046 169218 532102
rect 169274 532046 169342 532102
rect 169398 532046 169494 532102
rect 168874 531978 169494 532046
rect 168874 531922 168970 531978
rect 169026 531922 169094 531978
rect 169150 531922 169218 531978
rect 169274 531922 169342 531978
rect 169398 531922 169494 531978
rect 168874 527750 169494 531922
rect 183154 597212 183774 598268
rect 183154 597156 183250 597212
rect 183306 597156 183374 597212
rect 183430 597156 183498 597212
rect 183554 597156 183622 597212
rect 183678 597156 183774 597212
rect 183154 597088 183774 597156
rect 183154 597032 183250 597088
rect 183306 597032 183374 597088
rect 183430 597032 183498 597088
rect 183554 597032 183622 597088
rect 183678 597032 183774 597088
rect 183154 596964 183774 597032
rect 183154 596908 183250 596964
rect 183306 596908 183374 596964
rect 183430 596908 183498 596964
rect 183554 596908 183622 596964
rect 183678 596908 183774 596964
rect 183154 596840 183774 596908
rect 183154 596784 183250 596840
rect 183306 596784 183374 596840
rect 183430 596784 183498 596840
rect 183554 596784 183622 596840
rect 183678 596784 183774 596840
rect 183154 580350 183774 596784
rect 183154 580294 183250 580350
rect 183306 580294 183374 580350
rect 183430 580294 183498 580350
rect 183554 580294 183622 580350
rect 183678 580294 183774 580350
rect 183154 580226 183774 580294
rect 183154 580170 183250 580226
rect 183306 580170 183374 580226
rect 183430 580170 183498 580226
rect 183554 580170 183622 580226
rect 183678 580170 183774 580226
rect 183154 580102 183774 580170
rect 183154 580046 183250 580102
rect 183306 580046 183374 580102
rect 183430 580046 183498 580102
rect 183554 580046 183622 580102
rect 183678 580046 183774 580102
rect 183154 579978 183774 580046
rect 183154 579922 183250 579978
rect 183306 579922 183374 579978
rect 183430 579922 183498 579978
rect 183554 579922 183622 579978
rect 183678 579922 183774 579978
rect 183154 562350 183774 579922
rect 183154 562294 183250 562350
rect 183306 562294 183374 562350
rect 183430 562294 183498 562350
rect 183554 562294 183622 562350
rect 183678 562294 183774 562350
rect 183154 562226 183774 562294
rect 183154 562170 183250 562226
rect 183306 562170 183374 562226
rect 183430 562170 183498 562226
rect 183554 562170 183622 562226
rect 183678 562170 183774 562226
rect 183154 562102 183774 562170
rect 183154 562046 183250 562102
rect 183306 562046 183374 562102
rect 183430 562046 183498 562102
rect 183554 562046 183622 562102
rect 183678 562046 183774 562102
rect 183154 561978 183774 562046
rect 183154 561922 183250 561978
rect 183306 561922 183374 561978
rect 183430 561922 183498 561978
rect 183554 561922 183622 561978
rect 183678 561922 183774 561978
rect 183154 544350 183774 561922
rect 183154 544294 183250 544350
rect 183306 544294 183374 544350
rect 183430 544294 183498 544350
rect 183554 544294 183622 544350
rect 183678 544294 183774 544350
rect 183154 544226 183774 544294
rect 183154 544170 183250 544226
rect 183306 544170 183374 544226
rect 183430 544170 183498 544226
rect 183554 544170 183622 544226
rect 183678 544170 183774 544226
rect 183154 544102 183774 544170
rect 183154 544046 183250 544102
rect 183306 544046 183374 544102
rect 183430 544046 183498 544102
rect 183554 544046 183622 544102
rect 183678 544046 183774 544102
rect 183154 543978 183774 544046
rect 183154 543922 183250 543978
rect 183306 543922 183374 543978
rect 183430 543922 183498 543978
rect 183554 543922 183622 543978
rect 183678 543922 183774 543978
rect 183154 527750 183774 543922
rect 186874 598172 187494 598268
rect 186874 598116 186970 598172
rect 187026 598116 187094 598172
rect 187150 598116 187218 598172
rect 187274 598116 187342 598172
rect 187398 598116 187494 598172
rect 186874 598048 187494 598116
rect 186874 597992 186970 598048
rect 187026 597992 187094 598048
rect 187150 597992 187218 598048
rect 187274 597992 187342 598048
rect 187398 597992 187494 598048
rect 186874 597924 187494 597992
rect 186874 597868 186970 597924
rect 187026 597868 187094 597924
rect 187150 597868 187218 597924
rect 187274 597868 187342 597924
rect 187398 597868 187494 597924
rect 186874 597800 187494 597868
rect 186874 597744 186970 597800
rect 187026 597744 187094 597800
rect 187150 597744 187218 597800
rect 187274 597744 187342 597800
rect 187398 597744 187494 597800
rect 186874 586350 187494 597744
rect 186874 586294 186970 586350
rect 187026 586294 187094 586350
rect 187150 586294 187218 586350
rect 187274 586294 187342 586350
rect 187398 586294 187494 586350
rect 186874 586226 187494 586294
rect 186874 586170 186970 586226
rect 187026 586170 187094 586226
rect 187150 586170 187218 586226
rect 187274 586170 187342 586226
rect 187398 586170 187494 586226
rect 186874 586102 187494 586170
rect 186874 586046 186970 586102
rect 187026 586046 187094 586102
rect 187150 586046 187218 586102
rect 187274 586046 187342 586102
rect 187398 586046 187494 586102
rect 186874 585978 187494 586046
rect 186874 585922 186970 585978
rect 187026 585922 187094 585978
rect 187150 585922 187218 585978
rect 187274 585922 187342 585978
rect 187398 585922 187494 585978
rect 186874 568350 187494 585922
rect 186874 568294 186970 568350
rect 187026 568294 187094 568350
rect 187150 568294 187218 568350
rect 187274 568294 187342 568350
rect 187398 568294 187494 568350
rect 186874 568226 187494 568294
rect 186874 568170 186970 568226
rect 187026 568170 187094 568226
rect 187150 568170 187218 568226
rect 187274 568170 187342 568226
rect 187398 568170 187494 568226
rect 186874 568102 187494 568170
rect 186874 568046 186970 568102
rect 187026 568046 187094 568102
rect 187150 568046 187218 568102
rect 187274 568046 187342 568102
rect 187398 568046 187494 568102
rect 186874 567978 187494 568046
rect 186874 567922 186970 567978
rect 187026 567922 187094 567978
rect 187150 567922 187218 567978
rect 187274 567922 187342 567978
rect 187398 567922 187494 567978
rect 186874 550350 187494 567922
rect 186874 550294 186970 550350
rect 187026 550294 187094 550350
rect 187150 550294 187218 550350
rect 187274 550294 187342 550350
rect 187398 550294 187494 550350
rect 186874 550226 187494 550294
rect 186874 550170 186970 550226
rect 187026 550170 187094 550226
rect 187150 550170 187218 550226
rect 187274 550170 187342 550226
rect 187398 550170 187494 550226
rect 186874 550102 187494 550170
rect 186874 550046 186970 550102
rect 187026 550046 187094 550102
rect 187150 550046 187218 550102
rect 187274 550046 187342 550102
rect 187398 550046 187494 550102
rect 186874 549978 187494 550046
rect 186874 549922 186970 549978
rect 187026 549922 187094 549978
rect 187150 549922 187218 549978
rect 187274 549922 187342 549978
rect 187398 549922 187494 549978
rect 186874 532350 187494 549922
rect 186874 532294 186970 532350
rect 187026 532294 187094 532350
rect 187150 532294 187218 532350
rect 187274 532294 187342 532350
rect 187398 532294 187494 532350
rect 186874 532226 187494 532294
rect 186874 532170 186970 532226
rect 187026 532170 187094 532226
rect 187150 532170 187218 532226
rect 187274 532170 187342 532226
rect 187398 532170 187494 532226
rect 186874 532102 187494 532170
rect 186874 532046 186970 532102
rect 187026 532046 187094 532102
rect 187150 532046 187218 532102
rect 187274 532046 187342 532102
rect 187398 532046 187494 532102
rect 186874 531978 187494 532046
rect 186874 531922 186970 531978
rect 187026 531922 187094 531978
rect 187150 531922 187218 531978
rect 187274 531922 187342 531978
rect 187398 531922 187494 531978
rect 186874 527750 187494 531922
rect 201154 597212 201774 598268
rect 201154 597156 201250 597212
rect 201306 597156 201374 597212
rect 201430 597156 201498 597212
rect 201554 597156 201622 597212
rect 201678 597156 201774 597212
rect 201154 597088 201774 597156
rect 201154 597032 201250 597088
rect 201306 597032 201374 597088
rect 201430 597032 201498 597088
rect 201554 597032 201622 597088
rect 201678 597032 201774 597088
rect 201154 596964 201774 597032
rect 201154 596908 201250 596964
rect 201306 596908 201374 596964
rect 201430 596908 201498 596964
rect 201554 596908 201622 596964
rect 201678 596908 201774 596964
rect 201154 596840 201774 596908
rect 201154 596784 201250 596840
rect 201306 596784 201374 596840
rect 201430 596784 201498 596840
rect 201554 596784 201622 596840
rect 201678 596784 201774 596840
rect 201154 580350 201774 596784
rect 201154 580294 201250 580350
rect 201306 580294 201374 580350
rect 201430 580294 201498 580350
rect 201554 580294 201622 580350
rect 201678 580294 201774 580350
rect 201154 580226 201774 580294
rect 201154 580170 201250 580226
rect 201306 580170 201374 580226
rect 201430 580170 201498 580226
rect 201554 580170 201622 580226
rect 201678 580170 201774 580226
rect 201154 580102 201774 580170
rect 201154 580046 201250 580102
rect 201306 580046 201374 580102
rect 201430 580046 201498 580102
rect 201554 580046 201622 580102
rect 201678 580046 201774 580102
rect 201154 579978 201774 580046
rect 201154 579922 201250 579978
rect 201306 579922 201374 579978
rect 201430 579922 201498 579978
rect 201554 579922 201622 579978
rect 201678 579922 201774 579978
rect 201154 562350 201774 579922
rect 201154 562294 201250 562350
rect 201306 562294 201374 562350
rect 201430 562294 201498 562350
rect 201554 562294 201622 562350
rect 201678 562294 201774 562350
rect 201154 562226 201774 562294
rect 201154 562170 201250 562226
rect 201306 562170 201374 562226
rect 201430 562170 201498 562226
rect 201554 562170 201622 562226
rect 201678 562170 201774 562226
rect 201154 562102 201774 562170
rect 201154 562046 201250 562102
rect 201306 562046 201374 562102
rect 201430 562046 201498 562102
rect 201554 562046 201622 562102
rect 201678 562046 201774 562102
rect 201154 561978 201774 562046
rect 201154 561922 201250 561978
rect 201306 561922 201374 561978
rect 201430 561922 201498 561978
rect 201554 561922 201622 561978
rect 201678 561922 201774 561978
rect 201154 544350 201774 561922
rect 201154 544294 201250 544350
rect 201306 544294 201374 544350
rect 201430 544294 201498 544350
rect 201554 544294 201622 544350
rect 201678 544294 201774 544350
rect 201154 544226 201774 544294
rect 201154 544170 201250 544226
rect 201306 544170 201374 544226
rect 201430 544170 201498 544226
rect 201554 544170 201622 544226
rect 201678 544170 201774 544226
rect 201154 544102 201774 544170
rect 201154 544046 201250 544102
rect 201306 544046 201374 544102
rect 201430 544046 201498 544102
rect 201554 544046 201622 544102
rect 201678 544046 201774 544102
rect 201154 543978 201774 544046
rect 201154 543922 201250 543978
rect 201306 543922 201374 543978
rect 201430 543922 201498 543978
rect 201554 543922 201622 543978
rect 201678 543922 201774 543978
rect 201154 527750 201774 543922
rect 204874 598172 205494 598268
rect 204874 598116 204970 598172
rect 205026 598116 205094 598172
rect 205150 598116 205218 598172
rect 205274 598116 205342 598172
rect 205398 598116 205494 598172
rect 204874 598048 205494 598116
rect 204874 597992 204970 598048
rect 205026 597992 205094 598048
rect 205150 597992 205218 598048
rect 205274 597992 205342 598048
rect 205398 597992 205494 598048
rect 204874 597924 205494 597992
rect 204874 597868 204970 597924
rect 205026 597868 205094 597924
rect 205150 597868 205218 597924
rect 205274 597868 205342 597924
rect 205398 597868 205494 597924
rect 204874 597800 205494 597868
rect 204874 597744 204970 597800
rect 205026 597744 205094 597800
rect 205150 597744 205218 597800
rect 205274 597744 205342 597800
rect 205398 597744 205494 597800
rect 204874 586350 205494 597744
rect 204874 586294 204970 586350
rect 205026 586294 205094 586350
rect 205150 586294 205218 586350
rect 205274 586294 205342 586350
rect 205398 586294 205494 586350
rect 204874 586226 205494 586294
rect 204874 586170 204970 586226
rect 205026 586170 205094 586226
rect 205150 586170 205218 586226
rect 205274 586170 205342 586226
rect 205398 586170 205494 586226
rect 204874 586102 205494 586170
rect 204874 586046 204970 586102
rect 205026 586046 205094 586102
rect 205150 586046 205218 586102
rect 205274 586046 205342 586102
rect 205398 586046 205494 586102
rect 204874 585978 205494 586046
rect 204874 585922 204970 585978
rect 205026 585922 205094 585978
rect 205150 585922 205218 585978
rect 205274 585922 205342 585978
rect 205398 585922 205494 585978
rect 204874 568350 205494 585922
rect 204874 568294 204970 568350
rect 205026 568294 205094 568350
rect 205150 568294 205218 568350
rect 205274 568294 205342 568350
rect 205398 568294 205494 568350
rect 204874 568226 205494 568294
rect 204874 568170 204970 568226
rect 205026 568170 205094 568226
rect 205150 568170 205218 568226
rect 205274 568170 205342 568226
rect 205398 568170 205494 568226
rect 204874 568102 205494 568170
rect 204874 568046 204970 568102
rect 205026 568046 205094 568102
rect 205150 568046 205218 568102
rect 205274 568046 205342 568102
rect 205398 568046 205494 568102
rect 204874 567978 205494 568046
rect 204874 567922 204970 567978
rect 205026 567922 205094 567978
rect 205150 567922 205218 567978
rect 205274 567922 205342 567978
rect 205398 567922 205494 567978
rect 204874 550350 205494 567922
rect 204874 550294 204970 550350
rect 205026 550294 205094 550350
rect 205150 550294 205218 550350
rect 205274 550294 205342 550350
rect 205398 550294 205494 550350
rect 204874 550226 205494 550294
rect 204874 550170 204970 550226
rect 205026 550170 205094 550226
rect 205150 550170 205218 550226
rect 205274 550170 205342 550226
rect 205398 550170 205494 550226
rect 204874 550102 205494 550170
rect 204874 550046 204970 550102
rect 205026 550046 205094 550102
rect 205150 550046 205218 550102
rect 205274 550046 205342 550102
rect 205398 550046 205494 550102
rect 204874 549978 205494 550046
rect 204874 549922 204970 549978
rect 205026 549922 205094 549978
rect 205150 549922 205218 549978
rect 205274 549922 205342 549978
rect 205398 549922 205494 549978
rect 204874 532350 205494 549922
rect 204874 532294 204970 532350
rect 205026 532294 205094 532350
rect 205150 532294 205218 532350
rect 205274 532294 205342 532350
rect 205398 532294 205494 532350
rect 204874 532226 205494 532294
rect 204874 532170 204970 532226
rect 205026 532170 205094 532226
rect 205150 532170 205218 532226
rect 205274 532170 205342 532226
rect 205398 532170 205494 532226
rect 204874 532102 205494 532170
rect 204874 532046 204970 532102
rect 205026 532046 205094 532102
rect 205150 532046 205218 532102
rect 205274 532046 205342 532102
rect 205398 532046 205494 532102
rect 204874 531978 205494 532046
rect 204874 531922 204970 531978
rect 205026 531922 205094 531978
rect 205150 531922 205218 531978
rect 205274 531922 205342 531978
rect 205398 531922 205494 531978
rect 204874 527750 205494 531922
rect 219154 597212 219774 598268
rect 219154 597156 219250 597212
rect 219306 597156 219374 597212
rect 219430 597156 219498 597212
rect 219554 597156 219622 597212
rect 219678 597156 219774 597212
rect 219154 597088 219774 597156
rect 219154 597032 219250 597088
rect 219306 597032 219374 597088
rect 219430 597032 219498 597088
rect 219554 597032 219622 597088
rect 219678 597032 219774 597088
rect 219154 596964 219774 597032
rect 219154 596908 219250 596964
rect 219306 596908 219374 596964
rect 219430 596908 219498 596964
rect 219554 596908 219622 596964
rect 219678 596908 219774 596964
rect 219154 596840 219774 596908
rect 219154 596784 219250 596840
rect 219306 596784 219374 596840
rect 219430 596784 219498 596840
rect 219554 596784 219622 596840
rect 219678 596784 219774 596840
rect 219154 580350 219774 596784
rect 219154 580294 219250 580350
rect 219306 580294 219374 580350
rect 219430 580294 219498 580350
rect 219554 580294 219622 580350
rect 219678 580294 219774 580350
rect 219154 580226 219774 580294
rect 219154 580170 219250 580226
rect 219306 580170 219374 580226
rect 219430 580170 219498 580226
rect 219554 580170 219622 580226
rect 219678 580170 219774 580226
rect 219154 580102 219774 580170
rect 219154 580046 219250 580102
rect 219306 580046 219374 580102
rect 219430 580046 219498 580102
rect 219554 580046 219622 580102
rect 219678 580046 219774 580102
rect 219154 579978 219774 580046
rect 219154 579922 219250 579978
rect 219306 579922 219374 579978
rect 219430 579922 219498 579978
rect 219554 579922 219622 579978
rect 219678 579922 219774 579978
rect 219154 562350 219774 579922
rect 219154 562294 219250 562350
rect 219306 562294 219374 562350
rect 219430 562294 219498 562350
rect 219554 562294 219622 562350
rect 219678 562294 219774 562350
rect 219154 562226 219774 562294
rect 219154 562170 219250 562226
rect 219306 562170 219374 562226
rect 219430 562170 219498 562226
rect 219554 562170 219622 562226
rect 219678 562170 219774 562226
rect 219154 562102 219774 562170
rect 219154 562046 219250 562102
rect 219306 562046 219374 562102
rect 219430 562046 219498 562102
rect 219554 562046 219622 562102
rect 219678 562046 219774 562102
rect 219154 561978 219774 562046
rect 219154 561922 219250 561978
rect 219306 561922 219374 561978
rect 219430 561922 219498 561978
rect 219554 561922 219622 561978
rect 219678 561922 219774 561978
rect 219154 544350 219774 561922
rect 219154 544294 219250 544350
rect 219306 544294 219374 544350
rect 219430 544294 219498 544350
rect 219554 544294 219622 544350
rect 219678 544294 219774 544350
rect 219154 544226 219774 544294
rect 219154 544170 219250 544226
rect 219306 544170 219374 544226
rect 219430 544170 219498 544226
rect 219554 544170 219622 544226
rect 219678 544170 219774 544226
rect 219154 544102 219774 544170
rect 219154 544046 219250 544102
rect 219306 544046 219374 544102
rect 219430 544046 219498 544102
rect 219554 544046 219622 544102
rect 219678 544046 219774 544102
rect 219154 543978 219774 544046
rect 219154 543922 219250 543978
rect 219306 543922 219374 543978
rect 219430 543922 219498 543978
rect 219554 543922 219622 543978
rect 219678 543922 219774 543978
rect 219154 527750 219774 543922
rect 222874 598172 223494 598268
rect 222874 598116 222970 598172
rect 223026 598116 223094 598172
rect 223150 598116 223218 598172
rect 223274 598116 223342 598172
rect 223398 598116 223494 598172
rect 222874 598048 223494 598116
rect 222874 597992 222970 598048
rect 223026 597992 223094 598048
rect 223150 597992 223218 598048
rect 223274 597992 223342 598048
rect 223398 597992 223494 598048
rect 222874 597924 223494 597992
rect 222874 597868 222970 597924
rect 223026 597868 223094 597924
rect 223150 597868 223218 597924
rect 223274 597868 223342 597924
rect 223398 597868 223494 597924
rect 222874 597800 223494 597868
rect 222874 597744 222970 597800
rect 223026 597744 223094 597800
rect 223150 597744 223218 597800
rect 223274 597744 223342 597800
rect 223398 597744 223494 597800
rect 222874 586350 223494 597744
rect 222874 586294 222970 586350
rect 223026 586294 223094 586350
rect 223150 586294 223218 586350
rect 223274 586294 223342 586350
rect 223398 586294 223494 586350
rect 222874 586226 223494 586294
rect 222874 586170 222970 586226
rect 223026 586170 223094 586226
rect 223150 586170 223218 586226
rect 223274 586170 223342 586226
rect 223398 586170 223494 586226
rect 222874 586102 223494 586170
rect 222874 586046 222970 586102
rect 223026 586046 223094 586102
rect 223150 586046 223218 586102
rect 223274 586046 223342 586102
rect 223398 586046 223494 586102
rect 222874 585978 223494 586046
rect 222874 585922 222970 585978
rect 223026 585922 223094 585978
rect 223150 585922 223218 585978
rect 223274 585922 223342 585978
rect 223398 585922 223494 585978
rect 222874 568350 223494 585922
rect 222874 568294 222970 568350
rect 223026 568294 223094 568350
rect 223150 568294 223218 568350
rect 223274 568294 223342 568350
rect 223398 568294 223494 568350
rect 222874 568226 223494 568294
rect 222874 568170 222970 568226
rect 223026 568170 223094 568226
rect 223150 568170 223218 568226
rect 223274 568170 223342 568226
rect 223398 568170 223494 568226
rect 222874 568102 223494 568170
rect 222874 568046 222970 568102
rect 223026 568046 223094 568102
rect 223150 568046 223218 568102
rect 223274 568046 223342 568102
rect 223398 568046 223494 568102
rect 222874 567978 223494 568046
rect 222874 567922 222970 567978
rect 223026 567922 223094 567978
rect 223150 567922 223218 567978
rect 223274 567922 223342 567978
rect 223398 567922 223494 567978
rect 222874 550350 223494 567922
rect 222874 550294 222970 550350
rect 223026 550294 223094 550350
rect 223150 550294 223218 550350
rect 223274 550294 223342 550350
rect 223398 550294 223494 550350
rect 222874 550226 223494 550294
rect 222874 550170 222970 550226
rect 223026 550170 223094 550226
rect 223150 550170 223218 550226
rect 223274 550170 223342 550226
rect 223398 550170 223494 550226
rect 222874 550102 223494 550170
rect 222874 550046 222970 550102
rect 223026 550046 223094 550102
rect 223150 550046 223218 550102
rect 223274 550046 223342 550102
rect 223398 550046 223494 550102
rect 222874 549978 223494 550046
rect 222874 549922 222970 549978
rect 223026 549922 223094 549978
rect 223150 549922 223218 549978
rect 223274 549922 223342 549978
rect 223398 549922 223494 549978
rect 222874 532350 223494 549922
rect 222874 532294 222970 532350
rect 223026 532294 223094 532350
rect 223150 532294 223218 532350
rect 223274 532294 223342 532350
rect 223398 532294 223494 532350
rect 222874 532226 223494 532294
rect 222874 532170 222970 532226
rect 223026 532170 223094 532226
rect 223150 532170 223218 532226
rect 223274 532170 223342 532226
rect 223398 532170 223494 532226
rect 222874 532102 223494 532170
rect 222874 532046 222970 532102
rect 223026 532046 223094 532102
rect 223150 532046 223218 532102
rect 223274 532046 223342 532102
rect 223398 532046 223494 532102
rect 222874 531978 223494 532046
rect 222874 531922 222970 531978
rect 223026 531922 223094 531978
rect 223150 531922 223218 531978
rect 223274 531922 223342 531978
rect 223398 531922 223494 531978
rect 222874 528388 223494 531922
rect 237154 597212 237774 598268
rect 237154 597156 237250 597212
rect 237306 597156 237374 597212
rect 237430 597156 237498 597212
rect 237554 597156 237622 597212
rect 237678 597156 237774 597212
rect 237154 597088 237774 597156
rect 237154 597032 237250 597088
rect 237306 597032 237374 597088
rect 237430 597032 237498 597088
rect 237554 597032 237622 597088
rect 237678 597032 237774 597088
rect 237154 596964 237774 597032
rect 237154 596908 237250 596964
rect 237306 596908 237374 596964
rect 237430 596908 237498 596964
rect 237554 596908 237622 596964
rect 237678 596908 237774 596964
rect 237154 596840 237774 596908
rect 237154 596784 237250 596840
rect 237306 596784 237374 596840
rect 237430 596784 237498 596840
rect 237554 596784 237622 596840
rect 237678 596784 237774 596840
rect 237154 580350 237774 596784
rect 237154 580294 237250 580350
rect 237306 580294 237374 580350
rect 237430 580294 237498 580350
rect 237554 580294 237622 580350
rect 237678 580294 237774 580350
rect 237154 580226 237774 580294
rect 237154 580170 237250 580226
rect 237306 580170 237374 580226
rect 237430 580170 237498 580226
rect 237554 580170 237622 580226
rect 237678 580170 237774 580226
rect 237154 580102 237774 580170
rect 237154 580046 237250 580102
rect 237306 580046 237374 580102
rect 237430 580046 237498 580102
rect 237554 580046 237622 580102
rect 237678 580046 237774 580102
rect 237154 579978 237774 580046
rect 237154 579922 237250 579978
rect 237306 579922 237374 579978
rect 237430 579922 237498 579978
rect 237554 579922 237622 579978
rect 237678 579922 237774 579978
rect 237154 562350 237774 579922
rect 237154 562294 237250 562350
rect 237306 562294 237374 562350
rect 237430 562294 237498 562350
rect 237554 562294 237622 562350
rect 237678 562294 237774 562350
rect 237154 562226 237774 562294
rect 237154 562170 237250 562226
rect 237306 562170 237374 562226
rect 237430 562170 237498 562226
rect 237554 562170 237622 562226
rect 237678 562170 237774 562226
rect 237154 562102 237774 562170
rect 237154 562046 237250 562102
rect 237306 562046 237374 562102
rect 237430 562046 237498 562102
rect 237554 562046 237622 562102
rect 237678 562046 237774 562102
rect 237154 561978 237774 562046
rect 237154 561922 237250 561978
rect 237306 561922 237374 561978
rect 237430 561922 237498 561978
rect 237554 561922 237622 561978
rect 237678 561922 237774 561978
rect 237154 544350 237774 561922
rect 237154 544294 237250 544350
rect 237306 544294 237374 544350
rect 237430 544294 237498 544350
rect 237554 544294 237622 544350
rect 237678 544294 237774 544350
rect 237154 544226 237774 544294
rect 237154 544170 237250 544226
rect 237306 544170 237374 544226
rect 237430 544170 237498 544226
rect 237554 544170 237622 544226
rect 237678 544170 237774 544226
rect 237154 544102 237774 544170
rect 237154 544046 237250 544102
rect 237306 544046 237374 544102
rect 237430 544046 237498 544102
rect 237554 544046 237622 544102
rect 237678 544046 237774 544102
rect 237154 543978 237774 544046
rect 237154 543922 237250 543978
rect 237306 543922 237374 543978
rect 237430 543922 237498 543978
rect 237554 543922 237622 543978
rect 237678 543922 237774 543978
rect 237154 527750 237774 543922
rect 240874 598172 241494 598268
rect 240874 598116 240970 598172
rect 241026 598116 241094 598172
rect 241150 598116 241218 598172
rect 241274 598116 241342 598172
rect 241398 598116 241494 598172
rect 240874 598048 241494 598116
rect 240874 597992 240970 598048
rect 241026 597992 241094 598048
rect 241150 597992 241218 598048
rect 241274 597992 241342 598048
rect 241398 597992 241494 598048
rect 240874 597924 241494 597992
rect 240874 597868 240970 597924
rect 241026 597868 241094 597924
rect 241150 597868 241218 597924
rect 241274 597868 241342 597924
rect 241398 597868 241494 597924
rect 240874 597800 241494 597868
rect 240874 597744 240970 597800
rect 241026 597744 241094 597800
rect 241150 597744 241218 597800
rect 241274 597744 241342 597800
rect 241398 597744 241494 597800
rect 240874 586350 241494 597744
rect 240874 586294 240970 586350
rect 241026 586294 241094 586350
rect 241150 586294 241218 586350
rect 241274 586294 241342 586350
rect 241398 586294 241494 586350
rect 240874 586226 241494 586294
rect 240874 586170 240970 586226
rect 241026 586170 241094 586226
rect 241150 586170 241218 586226
rect 241274 586170 241342 586226
rect 241398 586170 241494 586226
rect 240874 586102 241494 586170
rect 240874 586046 240970 586102
rect 241026 586046 241094 586102
rect 241150 586046 241218 586102
rect 241274 586046 241342 586102
rect 241398 586046 241494 586102
rect 240874 585978 241494 586046
rect 240874 585922 240970 585978
rect 241026 585922 241094 585978
rect 241150 585922 241218 585978
rect 241274 585922 241342 585978
rect 241398 585922 241494 585978
rect 240874 568350 241494 585922
rect 240874 568294 240970 568350
rect 241026 568294 241094 568350
rect 241150 568294 241218 568350
rect 241274 568294 241342 568350
rect 241398 568294 241494 568350
rect 240874 568226 241494 568294
rect 240874 568170 240970 568226
rect 241026 568170 241094 568226
rect 241150 568170 241218 568226
rect 241274 568170 241342 568226
rect 241398 568170 241494 568226
rect 240874 568102 241494 568170
rect 240874 568046 240970 568102
rect 241026 568046 241094 568102
rect 241150 568046 241218 568102
rect 241274 568046 241342 568102
rect 241398 568046 241494 568102
rect 240874 567978 241494 568046
rect 240874 567922 240970 567978
rect 241026 567922 241094 567978
rect 241150 567922 241218 567978
rect 241274 567922 241342 567978
rect 241398 567922 241494 567978
rect 240874 550350 241494 567922
rect 240874 550294 240970 550350
rect 241026 550294 241094 550350
rect 241150 550294 241218 550350
rect 241274 550294 241342 550350
rect 241398 550294 241494 550350
rect 240874 550226 241494 550294
rect 240874 550170 240970 550226
rect 241026 550170 241094 550226
rect 241150 550170 241218 550226
rect 241274 550170 241342 550226
rect 241398 550170 241494 550226
rect 240874 550102 241494 550170
rect 240874 550046 240970 550102
rect 241026 550046 241094 550102
rect 241150 550046 241218 550102
rect 241274 550046 241342 550102
rect 241398 550046 241494 550102
rect 240874 549978 241494 550046
rect 240874 549922 240970 549978
rect 241026 549922 241094 549978
rect 241150 549922 241218 549978
rect 241274 549922 241342 549978
rect 241398 549922 241494 549978
rect 240874 532350 241494 549922
rect 240874 532294 240970 532350
rect 241026 532294 241094 532350
rect 241150 532294 241218 532350
rect 241274 532294 241342 532350
rect 241398 532294 241494 532350
rect 240874 532226 241494 532294
rect 240874 532170 240970 532226
rect 241026 532170 241094 532226
rect 241150 532170 241218 532226
rect 241274 532170 241342 532226
rect 241398 532170 241494 532226
rect 240874 532102 241494 532170
rect 240874 532046 240970 532102
rect 241026 532046 241094 532102
rect 241150 532046 241218 532102
rect 241274 532046 241342 532102
rect 241398 532046 241494 532102
rect 240874 531978 241494 532046
rect 240874 531922 240970 531978
rect 241026 531922 241094 531978
rect 241150 531922 241218 531978
rect 241274 531922 241342 531978
rect 241398 531922 241494 531978
rect 240874 527750 241494 531922
rect 255154 597212 255774 598268
rect 255154 597156 255250 597212
rect 255306 597156 255374 597212
rect 255430 597156 255498 597212
rect 255554 597156 255622 597212
rect 255678 597156 255774 597212
rect 255154 597088 255774 597156
rect 255154 597032 255250 597088
rect 255306 597032 255374 597088
rect 255430 597032 255498 597088
rect 255554 597032 255622 597088
rect 255678 597032 255774 597088
rect 255154 596964 255774 597032
rect 255154 596908 255250 596964
rect 255306 596908 255374 596964
rect 255430 596908 255498 596964
rect 255554 596908 255622 596964
rect 255678 596908 255774 596964
rect 255154 596840 255774 596908
rect 255154 596784 255250 596840
rect 255306 596784 255374 596840
rect 255430 596784 255498 596840
rect 255554 596784 255622 596840
rect 255678 596784 255774 596840
rect 255154 580350 255774 596784
rect 255154 580294 255250 580350
rect 255306 580294 255374 580350
rect 255430 580294 255498 580350
rect 255554 580294 255622 580350
rect 255678 580294 255774 580350
rect 255154 580226 255774 580294
rect 255154 580170 255250 580226
rect 255306 580170 255374 580226
rect 255430 580170 255498 580226
rect 255554 580170 255622 580226
rect 255678 580170 255774 580226
rect 255154 580102 255774 580170
rect 255154 580046 255250 580102
rect 255306 580046 255374 580102
rect 255430 580046 255498 580102
rect 255554 580046 255622 580102
rect 255678 580046 255774 580102
rect 255154 579978 255774 580046
rect 255154 579922 255250 579978
rect 255306 579922 255374 579978
rect 255430 579922 255498 579978
rect 255554 579922 255622 579978
rect 255678 579922 255774 579978
rect 255154 562350 255774 579922
rect 255154 562294 255250 562350
rect 255306 562294 255374 562350
rect 255430 562294 255498 562350
rect 255554 562294 255622 562350
rect 255678 562294 255774 562350
rect 255154 562226 255774 562294
rect 255154 562170 255250 562226
rect 255306 562170 255374 562226
rect 255430 562170 255498 562226
rect 255554 562170 255622 562226
rect 255678 562170 255774 562226
rect 255154 562102 255774 562170
rect 255154 562046 255250 562102
rect 255306 562046 255374 562102
rect 255430 562046 255498 562102
rect 255554 562046 255622 562102
rect 255678 562046 255774 562102
rect 255154 561978 255774 562046
rect 255154 561922 255250 561978
rect 255306 561922 255374 561978
rect 255430 561922 255498 561978
rect 255554 561922 255622 561978
rect 255678 561922 255774 561978
rect 255154 544350 255774 561922
rect 255154 544294 255250 544350
rect 255306 544294 255374 544350
rect 255430 544294 255498 544350
rect 255554 544294 255622 544350
rect 255678 544294 255774 544350
rect 255154 544226 255774 544294
rect 255154 544170 255250 544226
rect 255306 544170 255374 544226
rect 255430 544170 255498 544226
rect 255554 544170 255622 544226
rect 255678 544170 255774 544226
rect 255154 544102 255774 544170
rect 255154 544046 255250 544102
rect 255306 544046 255374 544102
rect 255430 544046 255498 544102
rect 255554 544046 255622 544102
rect 255678 544046 255774 544102
rect 255154 543978 255774 544046
rect 255154 543922 255250 543978
rect 255306 543922 255374 543978
rect 255430 543922 255498 543978
rect 255554 543922 255622 543978
rect 255678 543922 255774 543978
rect 255154 527750 255774 543922
rect 258874 598172 259494 598268
rect 258874 598116 258970 598172
rect 259026 598116 259094 598172
rect 259150 598116 259218 598172
rect 259274 598116 259342 598172
rect 259398 598116 259494 598172
rect 258874 598048 259494 598116
rect 258874 597992 258970 598048
rect 259026 597992 259094 598048
rect 259150 597992 259218 598048
rect 259274 597992 259342 598048
rect 259398 597992 259494 598048
rect 258874 597924 259494 597992
rect 258874 597868 258970 597924
rect 259026 597868 259094 597924
rect 259150 597868 259218 597924
rect 259274 597868 259342 597924
rect 259398 597868 259494 597924
rect 258874 597800 259494 597868
rect 258874 597744 258970 597800
rect 259026 597744 259094 597800
rect 259150 597744 259218 597800
rect 259274 597744 259342 597800
rect 259398 597744 259494 597800
rect 258874 586350 259494 597744
rect 258874 586294 258970 586350
rect 259026 586294 259094 586350
rect 259150 586294 259218 586350
rect 259274 586294 259342 586350
rect 259398 586294 259494 586350
rect 258874 586226 259494 586294
rect 258874 586170 258970 586226
rect 259026 586170 259094 586226
rect 259150 586170 259218 586226
rect 259274 586170 259342 586226
rect 259398 586170 259494 586226
rect 258874 586102 259494 586170
rect 258874 586046 258970 586102
rect 259026 586046 259094 586102
rect 259150 586046 259218 586102
rect 259274 586046 259342 586102
rect 259398 586046 259494 586102
rect 258874 585978 259494 586046
rect 258874 585922 258970 585978
rect 259026 585922 259094 585978
rect 259150 585922 259218 585978
rect 259274 585922 259342 585978
rect 259398 585922 259494 585978
rect 258874 568350 259494 585922
rect 258874 568294 258970 568350
rect 259026 568294 259094 568350
rect 259150 568294 259218 568350
rect 259274 568294 259342 568350
rect 259398 568294 259494 568350
rect 258874 568226 259494 568294
rect 258874 568170 258970 568226
rect 259026 568170 259094 568226
rect 259150 568170 259218 568226
rect 259274 568170 259342 568226
rect 259398 568170 259494 568226
rect 258874 568102 259494 568170
rect 258874 568046 258970 568102
rect 259026 568046 259094 568102
rect 259150 568046 259218 568102
rect 259274 568046 259342 568102
rect 259398 568046 259494 568102
rect 258874 567978 259494 568046
rect 258874 567922 258970 567978
rect 259026 567922 259094 567978
rect 259150 567922 259218 567978
rect 259274 567922 259342 567978
rect 259398 567922 259494 567978
rect 258874 550350 259494 567922
rect 258874 550294 258970 550350
rect 259026 550294 259094 550350
rect 259150 550294 259218 550350
rect 259274 550294 259342 550350
rect 259398 550294 259494 550350
rect 258874 550226 259494 550294
rect 258874 550170 258970 550226
rect 259026 550170 259094 550226
rect 259150 550170 259218 550226
rect 259274 550170 259342 550226
rect 259398 550170 259494 550226
rect 258874 550102 259494 550170
rect 258874 550046 258970 550102
rect 259026 550046 259094 550102
rect 259150 550046 259218 550102
rect 259274 550046 259342 550102
rect 259398 550046 259494 550102
rect 258874 549978 259494 550046
rect 258874 549922 258970 549978
rect 259026 549922 259094 549978
rect 259150 549922 259218 549978
rect 259274 549922 259342 549978
rect 259398 549922 259494 549978
rect 258874 532350 259494 549922
rect 258874 532294 258970 532350
rect 259026 532294 259094 532350
rect 259150 532294 259218 532350
rect 259274 532294 259342 532350
rect 259398 532294 259494 532350
rect 258874 532226 259494 532294
rect 258874 532170 258970 532226
rect 259026 532170 259094 532226
rect 259150 532170 259218 532226
rect 259274 532170 259342 532226
rect 259398 532170 259494 532226
rect 258874 532102 259494 532170
rect 258874 532046 258970 532102
rect 259026 532046 259094 532102
rect 259150 532046 259218 532102
rect 259274 532046 259342 532102
rect 259398 532046 259494 532102
rect 258874 531978 259494 532046
rect 258874 531922 258970 531978
rect 259026 531922 259094 531978
rect 259150 531922 259218 531978
rect 259274 531922 259342 531978
rect 259398 531922 259494 531978
rect 258874 527750 259494 531922
rect 273154 597212 273774 598268
rect 273154 597156 273250 597212
rect 273306 597156 273374 597212
rect 273430 597156 273498 597212
rect 273554 597156 273622 597212
rect 273678 597156 273774 597212
rect 273154 597088 273774 597156
rect 273154 597032 273250 597088
rect 273306 597032 273374 597088
rect 273430 597032 273498 597088
rect 273554 597032 273622 597088
rect 273678 597032 273774 597088
rect 273154 596964 273774 597032
rect 273154 596908 273250 596964
rect 273306 596908 273374 596964
rect 273430 596908 273498 596964
rect 273554 596908 273622 596964
rect 273678 596908 273774 596964
rect 273154 596840 273774 596908
rect 273154 596784 273250 596840
rect 273306 596784 273374 596840
rect 273430 596784 273498 596840
rect 273554 596784 273622 596840
rect 273678 596784 273774 596840
rect 273154 580350 273774 596784
rect 273154 580294 273250 580350
rect 273306 580294 273374 580350
rect 273430 580294 273498 580350
rect 273554 580294 273622 580350
rect 273678 580294 273774 580350
rect 273154 580226 273774 580294
rect 273154 580170 273250 580226
rect 273306 580170 273374 580226
rect 273430 580170 273498 580226
rect 273554 580170 273622 580226
rect 273678 580170 273774 580226
rect 273154 580102 273774 580170
rect 273154 580046 273250 580102
rect 273306 580046 273374 580102
rect 273430 580046 273498 580102
rect 273554 580046 273622 580102
rect 273678 580046 273774 580102
rect 273154 579978 273774 580046
rect 273154 579922 273250 579978
rect 273306 579922 273374 579978
rect 273430 579922 273498 579978
rect 273554 579922 273622 579978
rect 273678 579922 273774 579978
rect 273154 562350 273774 579922
rect 273154 562294 273250 562350
rect 273306 562294 273374 562350
rect 273430 562294 273498 562350
rect 273554 562294 273622 562350
rect 273678 562294 273774 562350
rect 273154 562226 273774 562294
rect 273154 562170 273250 562226
rect 273306 562170 273374 562226
rect 273430 562170 273498 562226
rect 273554 562170 273622 562226
rect 273678 562170 273774 562226
rect 273154 562102 273774 562170
rect 273154 562046 273250 562102
rect 273306 562046 273374 562102
rect 273430 562046 273498 562102
rect 273554 562046 273622 562102
rect 273678 562046 273774 562102
rect 273154 561978 273774 562046
rect 273154 561922 273250 561978
rect 273306 561922 273374 561978
rect 273430 561922 273498 561978
rect 273554 561922 273622 561978
rect 273678 561922 273774 561978
rect 273154 544350 273774 561922
rect 273154 544294 273250 544350
rect 273306 544294 273374 544350
rect 273430 544294 273498 544350
rect 273554 544294 273622 544350
rect 273678 544294 273774 544350
rect 273154 544226 273774 544294
rect 273154 544170 273250 544226
rect 273306 544170 273374 544226
rect 273430 544170 273498 544226
rect 273554 544170 273622 544226
rect 273678 544170 273774 544226
rect 273154 544102 273774 544170
rect 273154 544046 273250 544102
rect 273306 544046 273374 544102
rect 273430 544046 273498 544102
rect 273554 544046 273622 544102
rect 273678 544046 273774 544102
rect 273154 543978 273774 544046
rect 273154 543922 273250 543978
rect 273306 543922 273374 543978
rect 273430 543922 273498 543978
rect 273554 543922 273622 543978
rect 273678 543922 273774 543978
rect 273154 527750 273774 543922
rect 276874 598172 277494 598268
rect 276874 598116 276970 598172
rect 277026 598116 277094 598172
rect 277150 598116 277218 598172
rect 277274 598116 277342 598172
rect 277398 598116 277494 598172
rect 276874 598048 277494 598116
rect 276874 597992 276970 598048
rect 277026 597992 277094 598048
rect 277150 597992 277218 598048
rect 277274 597992 277342 598048
rect 277398 597992 277494 598048
rect 276874 597924 277494 597992
rect 276874 597868 276970 597924
rect 277026 597868 277094 597924
rect 277150 597868 277218 597924
rect 277274 597868 277342 597924
rect 277398 597868 277494 597924
rect 276874 597800 277494 597868
rect 276874 597744 276970 597800
rect 277026 597744 277094 597800
rect 277150 597744 277218 597800
rect 277274 597744 277342 597800
rect 277398 597744 277494 597800
rect 276874 586350 277494 597744
rect 276874 586294 276970 586350
rect 277026 586294 277094 586350
rect 277150 586294 277218 586350
rect 277274 586294 277342 586350
rect 277398 586294 277494 586350
rect 276874 586226 277494 586294
rect 276874 586170 276970 586226
rect 277026 586170 277094 586226
rect 277150 586170 277218 586226
rect 277274 586170 277342 586226
rect 277398 586170 277494 586226
rect 276874 586102 277494 586170
rect 276874 586046 276970 586102
rect 277026 586046 277094 586102
rect 277150 586046 277218 586102
rect 277274 586046 277342 586102
rect 277398 586046 277494 586102
rect 276874 585978 277494 586046
rect 276874 585922 276970 585978
rect 277026 585922 277094 585978
rect 277150 585922 277218 585978
rect 277274 585922 277342 585978
rect 277398 585922 277494 585978
rect 276874 568350 277494 585922
rect 276874 568294 276970 568350
rect 277026 568294 277094 568350
rect 277150 568294 277218 568350
rect 277274 568294 277342 568350
rect 277398 568294 277494 568350
rect 276874 568226 277494 568294
rect 276874 568170 276970 568226
rect 277026 568170 277094 568226
rect 277150 568170 277218 568226
rect 277274 568170 277342 568226
rect 277398 568170 277494 568226
rect 276874 568102 277494 568170
rect 276874 568046 276970 568102
rect 277026 568046 277094 568102
rect 277150 568046 277218 568102
rect 277274 568046 277342 568102
rect 277398 568046 277494 568102
rect 276874 567978 277494 568046
rect 276874 567922 276970 567978
rect 277026 567922 277094 567978
rect 277150 567922 277218 567978
rect 277274 567922 277342 567978
rect 277398 567922 277494 567978
rect 276874 550350 277494 567922
rect 276874 550294 276970 550350
rect 277026 550294 277094 550350
rect 277150 550294 277218 550350
rect 277274 550294 277342 550350
rect 277398 550294 277494 550350
rect 276874 550226 277494 550294
rect 276874 550170 276970 550226
rect 277026 550170 277094 550226
rect 277150 550170 277218 550226
rect 277274 550170 277342 550226
rect 277398 550170 277494 550226
rect 276874 550102 277494 550170
rect 276874 550046 276970 550102
rect 277026 550046 277094 550102
rect 277150 550046 277218 550102
rect 277274 550046 277342 550102
rect 277398 550046 277494 550102
rect 276874 549978 277494 550046
rect 276874 549922 276970 549978
rect 277026 549922 277094 549978
rect 277150 549922 277218 549978
rect 277274 549922 277342 549978
rect 277398 549922 277494 549978
rect 276874 532350 277494 549922
rect 276874 532294 276970 532350
rect 277026 532294 277094 532350
rect 277150 532294 277218 532350
rect 277274 532294 277342 532350
rect 277398 532294 277494 532350
rect 276874 532226 277494 532294
rect 276874 532170 276970 532226
rect 277026 532170 277094 532226
rect 277150 532170 277218 532226
rect 277274 532170 277342 532226
rect 277398 532170 277494 532226
rect 276874 532102 277494 532170
rect 276874 532046 276970 532102
rect 277026 532046 277094 532102
rect 277150 532046 277218 532102
rect 277274 532046 277342 532102
rect 277398 532046 277494 532102
rect 276874 531978 277494 532046
rect 276874 531922 276970 531978
rect 277026 531922 277094 531978
rect 277150 531922 277218 531978
rect 277274 531922 277342 531978
rect 277398 531922 277494 531978
rect 276874 527750 277494 531922
rect 291154 597212 291774 598268
rect 291154 597156 291250 597212
rect 291306 597156 291374 597212
rect 291430 597156 291498 597212
rect 291554 597156 291622 597212
rect 291678 597156 291774 597212
rect 291154 597088 291774 597156
rect 291154 597032 291250 597088
rect 291306 597032 291374 597088
rect 291430 597032 291498 597088
rect 291554 597032 291622 597088
rect 291678 597032 291774 597088
rect 291154 596964 291774 597032
rect 291154 596908 291250 596964
rect 291306 596908 291374 596964
rect 291430 596908 291498 596964
rect 291554 596908 291622 596964
rect 291678 596908 291774 596964
rect 291154 596840 291774 596908
rect 291154 596784 291250 596840
rect 291306 596784 291374 596840
rect 291430 596784 291498 596840
rect 291554 596784 291622 596840
rect 291678 596784 291774 596840
rect 291154 580350 291774 596784
rect 291154 580294 291250 580350
rect 291306 580294 291374 580350
rect 291430 580294 291498 580350
rect 291554 580294 291622 580350
rect 291678 580294 291774 580350
rect 291154 580226 291774 580294
rect 291154 580170 291250 580226
rect 291306 580170 291374 580226
rect 291430 580170 291498 580226
rect 291554 580170 291622 580226
rect 291678 580170 291774 580226
rect 291154 580102 291774 580170
rect 291154 580046 291250 580102
rect 291306 580046 291374 580102
rect 291430 580046 291498 580102
rect 291554 580046 291622 580102
rect 291678 580046 291774 580102
rect 291154 579978 291774 580046
rect 291154 579922 291250 579978
rect 291306 579922 291374 579978
rect 291430 579922 291498 579978
rect 291554 579922 291622 579978
rect 291678 579922 291774 579978
rect 291154 562350 291774 579922
rect 291154 562294 291250 562350
rect 291306 562294 291374 562350
rect 291430 562294 291498 562350
rect 291554 562294 291622 562350
rect 291678 562294 291774 562350
rect 291154 562226 291774 562294
rect 291154 562170 291250 562226
rect 291306 562170 291374 562226
rect 291430 562170 291498 562226
rect 291554 562170 291622 562226
rect 291678 562170 291774 562226
rect 291154 562102 291774 562170
rect 291154 562046 291250 562102
rect 291306 562046 291374 562102
rect 291430 562046 291498 562102
rect 291554 562046 291622 562102
rect 291678 562046 291774 562102
rect 291154 561978 291774 562046
rect 291154 561922 291250 561978
rect 291306 561922 291374 561978
rect 291430 561922 291498 561978
rect 291554 561922 291622 561978
rect 291678 561922 291774 561978
rect 291154 544350 291774 561922
rect 291154 544294 291250 544350
rect 291306 544294 291374 544350
rect 291430 544294 291498 544350
rect 291554 544294 291622 544350
rect 291678 544294 291774 544350
rect 291154 544226 291774 544294
rect 291154 544170 291250 544226
rect 291306 544170 291374 544226
rect 291430 544170 291498 544226
rect 291554 544170 291622 544226
rect 291678 544170 291774 544226
rect 291154 544102 291774 544170
rect 291154 544046 291250 544102
rect 291306 544046 291374 544102
rect 291430 544046 291498 544102
rect 291554 544046 291622 544102
rect 291678 544046 291774 544102
rect 291154 543978 291774 544046
rect 291154 543922 291250 543978
rect 291306 543922 291374 543978
rect 291430 543922 291498 543978
rect 291554 543922 291622 543978
rect 291678 543922 291774 543978
rect 291154 527750 291774 543922
rect 294874 598172 295494 598268
rect 294874 598116 294970 598172
rect 295026 598116 295094 598172
rect 295150 598116 295218 598172
rect 295274 598116 295342 598172
rect 295398 598116 295494 598172
rect 294874 598048 295494 598116
rect 294874 597992 294970 598048
rect 295026 597992 295094 598048
rect 295150 597992 295218 598048
rect 295274 597992 295342 598048
rect 295398 597992 295494 598048
rect 294874 597924 295494 597992
rect 294874 597868 294970 597924
rect 295026 597868 295094 597924
rect 295150 597868 295218 597924
rect 295274 597868 295342 597924
rect 295398 597868 295494 597924
rect 294874 597800 295494 597868
rect 294874 597744 294970 597800
rect 295026 597744 295094 597800
rect 295150 597744 295218 597800
rect 295274 597744 295342 597800
rect 295398 597744 295494 597800
rect 294874 586350 295494 597744
rect 294874 586294 294970 586350
rect 295026 586294 295094 586350
rect 295150 586294 295218 586350
rect 295274 586294 295342 586350
rect 295398 586294 295494 586350
rect 294874 586226 295494 586294
rect 294874 586170 294970 586226
rect 295026 586170 295094 586226
rect 295150 586170 295218 586226
rect 295274 586170 295342 586226
rect 295398 586170 295494 586226
rect 294874 586102 295494 586170
rect 294874 586046 294970 586102
rect 295026 586046 295094 586102
rect 295150 586046 295218 586102
rect 295274 586046 295342 586102
rect 295398 586046 295494 586102
rect 294874 585978 295494 586046
rect 294874 585922 294970 585978
rect 295026 585922 295094 585978
rect 295150 585922 295218 585978
rect 295274 585922 295342 585978
rect 295398 585922 295494 585978
rect 294874 568350 295494 585922
rect 294874 568294 294970 568350
rect 295026 568294 295094 568350
rect 295150 568294 295218 568350
rect 295274 568294 295342 568350
rect 295398 568294 295494 568350
rect 294874 568226 295494 568294
rect 294874 568170 294970 568226
rect 295026 568170 295094 568226
rect 295150 568170 295218 568226
rect 295274 568170 295342 568226
rect 295398 568170 295494 568226
rect 294874 568102 295494 568170
rect 294874 568046 294970 568102
rect 295026 568046 295094 568102
rect 295150 568046 295218 568102
rect 295274 568046 295342 568102
rect 295398 568046 295494 568102
rect 294874 567978 295494 568046
rect 294874 567922 294970 567978
rect 295026 567922 295094 567978
rect 295150 567922 295218 567978
rect 295274 567922 295342 567978
rect 295398 567922 295494 567978
rect 294874 550350 295494 567922
rect 294874 550294 294970 550350
rect 295026 550294 295094 550350
rect 295150 550294 295218 550350
rect 295274 550294 295342 550350
rect 295398 550294 295494 550350
rect 294874 550226 295494 550294
rect 294874 550170 294970 550226
rect 295026 550170 295094 550226
rect 295150 550170 295218 550226
rect 295274 550170 295342 550226
rect 295398 550170 295494 550226
rect 294874 550102 295494 550170
rect 294874 550046 294970 550102
rect 295026 550046 295094 550102
rect 295150 550046 295218 550102
rect 295274 550046 295342 550102
rect 295398 550046 295494 550102
rect 294874 549978 295494 550046
rect 294874 549922 294970 549978
rect 295026 549922 295094 549978
rect 295150 549922 295218 549978
rect 295274 549922 295342 549978
rect 295398 549922 295494 549978
rect 294874 532350 295494 549922
rect 294874 532294 294970 532350
rect 295026 532294 295094 532350
rect 295150 532294 295218 532350
rect 295274 532294 295342 532350
rect 295398 532294 295494 532350
rect 294874 532226 295494 532294
rect 294874 532170 294970 532226
rect 295026 532170 295094 532226
rect 295150 532170 295218 532226
rect 295274 532170 295342 532226
rect 295398 532170 295494 532226
rect 294874 532102 295494 532170
rect 294874 532046 294970 532102
rect 295026 532046 295094 532102
rect 295150 532046 295218 532102
rect 295274 532046 295342 532102
rect 295398 532046 295494 532102
rect 294874 531978 295494 532046
rect 294874 531922 294970 531978
rect 295026 531922 295094 531978
rect 295150 531922 295218 531978
rect 295274 531922 295342 531978
rect 295398 531922 295494 531978
rect 294874 527750 295494 531922
rect 309154 597212 309774 598268
rect 309154 597156 309250 597212
rect 309306 597156 309374 597212
rect 309430 597156 309498 597212
rect 309554 597156 309622 597212
rect 309678 597156 309774 597212
rect 309154 597088 309774 597156
rect 309154 597032 309250 597088
rect 309306 597032 309374 597088
rect 309430 597032 309498 597088
rect 309554 597032 309622 597088
rect 309678 597032 309774 597088
rect 309154 596964 309774 597032
rect 309154 596908 309250 596964
rect 309306 596908 309374 596964
rect 309430 596908 309498 596964
rect 309554 596908 309622 596964
rect 309678 596908 309774 596964
rect 309154 596840 309774 596908
rect 309154 596784 309250 596840
rect 309306 596784 309374 596840
rect 309430 596784 309498 596840
rect 309554 596784 309622 596840
rect 309678 596784 309774 596840
rect 309154 580350 309774 596784
rect 309154 580294 309250 580350
rect 309306 580294 309374 580350
rect 309430 580294 309498 580350
rect 309554 580294 309622 580350
rect 309678 580294 309774 580350
rect 309154 580226 309774 580294
rect 309154 580170 309250 580226
rect 309306 580170 309374 580226
rect 309430 580170 309498 580226
rect 309554 580170 309622 580226
rect 309678 580170 309774 580226
rect 309154 580102 309774 580170
rect 309154 580046 309250 580102
rect 309306 580046 309374 580102
rect 309430 580046 309498 580102
rect 309554 580046 309622 580102
rect 309678 580046 309774 580102
rect 309154 579978 309774 580046
rect 309154 579922 309250 579978
rect 309306 579922 309374 579978
rect 309430 579922 309498 579978
rect 309554 579922 309622 579978
rect 309678 579922 309774 579978
rect 309154 562350 309774 579922
rect 309154 562294 309250 562350
rect 309306 562294 309374 562350
rect 309430 562294 309498 562350
rect 309554 562294 309622 562350
rect 309678 562294 309774 562350
rect 309154 562226 309774 562294
rect 309154 562170 309250 562226
rect 309306 562170 309374 562226
rect 309430 562170 309498 562226
rect 309554 562170 309622 562226
rect 309678 562170 309774 562226
rect 309154 562102 309774 562170
rect 309154 562046 309250 562102
rect 309306 562046 309374 562102
rect 309430 562046 309498 562102
rect 309554 562046 309622 562102
rect 309678 562046 309774 562102
rect 309154 561978 309774 562046
rect 309154 561922 309250 561978
rect 309306 561922 309374 561978
rect 309430 561922 309498 561978
rect 309554 561922 309622 561978
rect 309678 561922 309774 561978
rect 309154 544350 309774 561922
rect 309154 544294 309250 544350
rect 309306 544294 309374 544350
rect 309430 544294 309498 544350
rect 309554 544294 309622 544350
rect 309678 544294 309774 544350
rect 309154 544226 309774 544294
rect 309154 544170 309250 544226
rect 309306 544170 309374 544226
rect 309430 544170 309498 544226
rect 309554 544170 309622 544226
rect 309678 544170 309774 544226
rect 309154 544102 309774 544170
rect 309154 544046 309250 544102
rect 309306 544046 309374 544102
rect 309430 544046 309498 544102
rect 309554 544046 309622 544102
rect 309678 544046 309774 544102
rect 309154 543978 309774 544046
rect 309154 543922 309250 543978
rect 309306 543922 309374 543978
rect 309430 543922 309498 543978
rect 309554 543922 309622 543978
rect 309678 543922 309774 543978
rect 309154 527750 309774 543922
rect 312874 598172 313494 598268
rect 312874 598116 312970 598172
rect 313026 598116 313094 598172
rect 313150 598116 313218 598172
rect 313274 598116 313342 598172
rect 313398 598116 313494 598172
rect 312874 598048 313494 598116
rect 312874 597992 312970 598048
rect 313026 597992 313094 598048
rect 313150 597992 313218 598048
rect 313274 597992 313342 598048
rect 313398 597992 313494 598048
rect 312874 597924 313494 597992
rect 312874 597868 312970 597924
rect 313026 597868 313094 597924
rect 313150 597868 313218 597924
rect 313274 597868 313342 597924
rect 313398 597868 313494 597924
rect 312874 597800 313494 597868
rect 312874 597744 312970 597800
rect 313026 597744 313094 597800
rect 313150 597744 313218 597800
rect 313274 597744 313342 597800
rect 313398 597744 313494 597800
rect 312874 586350 313494 597744
rect 312874 586294 312970 586350
rect 313026 586294 313094 586350
rect 313150 586294 313218 586350
rect 313274 586294 313342 586350
rect 313398 586294 313494 586350
rect 312874 586226 313494 586294
rect 312874 586170 312970 586226
rect 313026 586170 313094 586226
rect 313150 586170 313218 586226
rect 313274 586170 313342 586226
rect 313398 586170 313494 586226
rect 312874 586102 313494 586170
rect 312874 586046 312970 586102
rect 313026 586046 313094 586102
rect 313150 586046 313218 586102
rect 313274 586046 313342 586102
rect 313398 586046 313494 586102
rect 312874 585978 313494 586046
rect 312874 585922 312970 585978
rect 313026 585922 313094 585978
rect 313150 585922 313218 585978
rect 313274 585922 313342 585978
rect 313398 585922 313494 585978
rect 312874 568350 313494 585922
rect 312874 568294 312970 568350
rect 313026 568294 313094 568350
rect 313150 568294 313218 568350
rect 313274 568294 313342 568350
rect 313398 568294 313494 568350
rect 312874 568226 313494 568294
rect 312874 568170 312970 568226
rect 313026 568170 313094 568226
rect 313150 568170 313218 568226
rect 313274 568170 313342 568226
rect 313398 568170 313494 568226
rect 312874 568102 313494 568170
rect 312874 568046 312970 568102
rect 313026 568046 313094 568102
rect 313150 568046 313218 568102
rect 313274 568046 313342 568102
rect 313398 568046 313494 568102
rect 312874 567978 313494 568046
rect 312874 567922 312970 567978
rect 313026 567922 313094 567978
rect 313150 567922 313218 567978
rect 313274 567922 313342 567978
rect 313398 567922 313494 567978
rect 312874 550350 313494 567922
rect 312874 550294 312970 550350
rect 313026 550294 313094 550350
rect 313150 550294 313218 550350
rect 313274 550294 313342 550350
rect 313398 550294 313494 550350
rect 312874 550226 313494 550294
rect 312874 550170 312970 550226
rect 313026 550170 313094 550226
rect 313150 550170 313218 550226
rect 313274 550170 313342 550226
rect 313398 550170 313494 550226
rect 312874 550102 313494 550170
rect 312874 550046 312970 550102
rect 313026 550046 313094 550102
rect 313150 550046 313218 550102
rect 313274 550046 313342 550102
rect 313398 550046 313494 550102
rect 312874 549978 313494 550046
rect 312874 549922 312970 549978
rect 313026 549922 313094 549978
rect 313150 549922 313218 549978
rect 313274 549922 313342 549978
rect 313398 549922 313494 549978
rect 312874 532350 313494 549922
rect 312874 532294 312970 532350
rect 313026 532294 313094 532350
rect 313150 532294 313218 532350
rect 313274 532294 313342 532350
rect 313398 532294 313494 532350
rect 312874 532226 313494 532294
rect 312874 532170 312970 532226
rect 313026 532170 313094 532226
rect 313150 532170 313218 532226
rect 313274 532170 313342 532226
rect 313398 532170 313494 532226
rect 312874 532102 313494 532170
rect 312874 532046 312970 532102
rect 313026 532046 313094 532102
rect 313150 532046 313218 532102
rect 313274 532046 313342 532102
rect 313398 532046 313494 532102
rect 312874 531978 313494 532046
rect 312874 531922 312970 531978
rect 313026 531922 313094 531978
rect 313150 531922 313218 531978
rect 313274 531922 313342 531978
rect 313398 531922 313494 531978
rect 312874 527750 313494 531922
rect 327154 597212 327774 598268
rect 327154 597156 327250 597212
rect 327306 597156 327374 597212
rect 327430 597156 327498 597212
rect 327554 597156 327622 597212
rect 327678 597156 327774 597212
rect 327154 597088 327774 597156
rect 327154 597032 327250 597088
rect 327306 597032 327374 597088
rect 327430 597032 327498 597088
rect 327554 597032 327622 597088
rect 327678 597032 327774 597088
rect 327154 596964 327774 597032
rect 327154 596908 327250 596964
rect 327306 596908 327374 596964
rect 327430 596908 327498 596964
rect 327554 596908 327622 596964
rect 327678 596908 327774 596964
rect 327154 596840 327774 596908
rect 327154 596784 327250 596840
rect 327306 596784 327374 596840
rect 327430 596784 327498 596840
rect 327554 596784 327622 596840
rect 327678 596784 327774 596840
rect 327154 580350 327774 596784
rect 327154 580294 327250 580350
rect 327306 580294 327374 580350
rect 327430 580294 327498 580350
rect 327554 580294 327622 580350
rect 327678 580294 327774 580350
rect 327154 580226 327774 580294
rect 327154 580170 327250 580226
rect 327306 580170 327374 580226
rect 327430 580170 327498 580226
rect 327554 580170 327622 580226
rect 327678 580170 327774 580226
rect 327154 580102 327774 580170
rect 327154 580046 327250 580102
rect 327306 580046 327374 580102
rect 327430 580046 327498 580102
rect 327554 580046 327622 580102
rect 327678 580046 327774 580102
rect 327154 579978 327774 580046
rect 327154 579922 327250 579978
rect 327306 579922 327374 579978
rect 327430 579922 327498 579978
rect 327554 579922 327622 579978
rect 327678 579922 327774 579978
rect 327154 562350 327774 579922
rect 327154 562294 327250 562350
rect 327306 562294 327374 562350
rect 327430 562294 327498 562350
rect 327554 562294 327622 562350
rect 327678 562294 327774 562350
rect 327154 562226 327774 562294
rect 327154 562170 327250 562226
rect 327306 562170 327374 562226
rect 327430 562170 327498 562226
rect 327554 562170 327622 562226
rect 327678 562170 327774 562226
rect 327154 562102 327774 562170
rect 327154 562046 327250 562102
rect 327306 562046 327374 562102
rect 327430 562046 327498 562102
rect 327554 562046 327622 562102
rect 327678 562046 327774 562102
rect 327154 561978 327774 562046
rect 327154 561922 327250 561978
rect 327306 561922 327374 561978
rect 327430 561922 327498 561978
rect 327554 561922 327622 561978
rect 327678 561922 327774 561978
rect 327154 544350 327774 561922
rect 327154 544294 327250 544350
rect 327306 544294 327374 544350
rect 327430 544294 327498 544350
rect 327554 544294 327622 544350
rect 327678 544294 327774 544350
rect 327154 544226 327774 544294
rect 327154 544170 327250 544226
rect 327306 544170 327374 544226
rect 327430 544170 327498 544226
rect 327554 544170 327622 544226
rect 327678 544170 327774 544226
rect 327154 544102 327774 544170
rect 327154 544046 327250 544102
rect 327306 544046 327374 544102
rect 327430 544046 327498 544102
rect 327554 544046 327622 544102
rect 327678 544046 327774 544102
rect 327154 543978 327774 544046
rect 327154 543922 327250 543978
rect 327306 543922 327374 543978
rect 327430 543922 327498 543978
rect 327554 543922 327622 543978
rect 327678 543922 327774 543978
rect 327154 527750 327774 543922
rect 330874 598172 331494 598268
rect 330874 598116 330970 598172
rect 331026 598116 331094 598172
rect 331150 598116 331218 598172
rect 331274 598116 331342 598172
rect 331398 598116 331494 598172
rect 330874 598048 331494 598116
rect 330874 597992 330970 598048
rect 331026 597992 331094 598048
rect 331150 597992 331218 598048
rect 331274 597992 331342 598048
rect 331398 597992 331494 598048
rect 330874 597924 331494 597992
rect 330874 597868 330970 597924
rect 331026 597868 331094 597924
rect 331150 597868 331218 597924
rect 331274 597868 331342 597924
rect 331398 597868 331494 597924
rect 330874 597800 331494 597868
rect 330874 597744 330970 597800
rect 331026 597744 331094 597800
rect 331150 597744 331218 597800
rect 331274 597744 331342 597800
rect 331398 597744 331494 597800
rect 330874 586350 331494 597744
rect 330874 586294 330970 586350
rect 331026 586294 331094 586350
rect 331150 586294 331218 586350
rect 331274 586294 331342 586350
rect 331398 586294 331494 586350
rect 330874 586226 331494 586294
rect 330874 586170 330970 586226
rect 331026 586170 331094 586226
rect 331150 586170 331218 586226
rect 331274 586170 331342 586226
rect 331398 586170 331494 586226
rect 330874 586102 331494 586170
rect 330874 586046 330970 586102
rect 331026 586046 331094 586102
rect 331150 586046 331218 586102
rect 331274 586046 331342 586102
rect 331398 586046 331494 586102
rect 330874 585978 331494 586046
rect 330874 585922 330970 585978
rect 331026 585922 331094 585978
rect 331150 585922 331218 585978
rect 331274 585922 331342 585978
rect 331398 585922 331494 585978
rect 330874 568350 331494 585922
rect 330874 568294 330970 568350
rect 331026 568294 331094 568350
rect 331150 568294 331218 568350
rect 331274 568294 331342 568350
rect 331398 568294 331494 568350
rect 330874 568226 331494 568294
rect 330874 568170 330970 568226
rect 331026 568170 331094 568226
rect 331150 568170 331218 568226
rect 331274 568170 331342 568226
rect 331398 568170 331494 568226
rect 330874 568102 331494 568170
rect 330874 568046 330970 568102
rect 331026 568046 331094 568102
rect 331150 568046 331218 568102
rect 331274 568046 331342 568102
rect 331398 568046 331494 568102
rect 330874 567978 331494 568046
rect 330874 567922 330970 567978
rect 331026 567922 331094 567978
rect 331150 567922 331218 567978
rect 331274 567922 331342 567978
rect 331398 567922 331494 567978
rect 330874 550350 331494 567922
rect 330874 550294 330970 550350
rect 331026 550294 331094 550350
rect 331150 550294 331218 550350
rect 331274 550294 331342 550350
rect 331398 550294 331494 550350
rect 330874 550226 331494 550294
rect 330874 550170 330970 550226
rect 331026 550170 331094 550226
rect 331150 550170 331218 550226
rect 331274 550170 331342 550226
rect 331398 550170 331494 550226
rect 330874 550102 331494 550170
rect 330874 550046 330970 550102
rect 331026 550046 331094 550102
rect 331150 550046 331218 550102
rect 331274 550046 331342 550102
rect 331398 550046 331494 550102
rect 330874 549978 331494 550046
rect 330874 549922 330970 549978
rect 331026 549922 331094 549978
rect 331150 549922 331218 549978
rect 331274 549922 331342 549978
rect 331398 549922 331494 549978
rect 330874 532350 331494 549922
rect 330874 532294 330970 532350
rect 331026 532294 331094 532350
rect 331150 532294 331218 532350
rect 331274 532294 331342 532350
rect 331398 532294 331494 532350
rect 330874 532226 331494 532294
rect 330874 532170 330970 532226
rect 331026 532170 331094 532226
rect 331150 532170 331218 532226
rect 331274 532170 331342 532226
rect 331398 532170 331494 532226
rect 330874 532102 331494 532170
rect 330874 532046 330970 532102
rect 331026 532046 331094 532102
rect 331150 532046 331218 532102
rect 331274 532046 331342 532102
rect 331398 532046 331494 532102
rect 330874 531978 331494 532046
rect 330874 531922 330970 531978
rect 331026 531922 331094 531978
rect 331150 531922 331218 531978
rect 331274 531922 331342 531978
rect 331398 531922 331494 531978
rect 330874 528388 331494 531922
rect 345154 597212 345774 598268
rect 345154 597156 345250 597212
rect 345306 597156 345374 597212
rect 345430 597156 345498 597212
rect 345554 597156 345622 597212
rect 345678 597156 345774 597212
rect 345154 597088 345774 597156
rect 345154 597032 345250 597088
rect 345306 597032 345374 597088
rect 345430 597032 345498 597088
rect 345554 597032 345622 597088
rect 345678 597032 345774 597088
rect 345154 596964 345774 597032
rect 345154 596908 345250 596964
rect 345306 596908 345374 596964
rect 345430 596908 345498 596964
rect 345554 596908 345622 596964
rect 345678 596908 345774 596964
rect 345154 596840 345774 596908
rect 345154 596784 345250 596840
rect 345306 596784 345374 596840
rect 345430 596784 345498 596840
rect 345554 596784 345622 596840
rect 345678 596784 345774 596840
rect 345154 580350 345774 596784
rect 345154 580294 345250 580350
rect 345306 580294 345374 580350
rect 345430 580294 345498 580350
rect 345554 580294 345622 580350
rect 345678 580294 345774 580350
rect 345154 580226 345774 580294
rect 345154 580170 345250 580226
rect 345306 580170 345374 580226
rect 345430 580170 345498 580226
rect 345554 580170 345622 580226
rect 345678 580170 345774 580226
rect 345154 580102 345774 580170
rect 345154 580046 345250 580102
rect 345306 580046 345374 580102
rect 345430 580046 345498 580102
rect 345554 580046 345622 580102
rect 345678 580046 345774 580102
rect 345154 579978 345774 580046
rect 345154 579922 345250 579978
rect 345306 579922 345374 579978
rect 345430 579922 345498 579978
rect 345554 579922 345622 579978
rect 345678 579922 345774 579978
rect 345154 562350 345774 579922
rect 345154 562294 345250 562350
rect 345306 562294 345374 562350
rect 345430 562294 345498 562350
rect 345554 562294 345622 562350
rect 345678 562294 345774 562350
rect 345154 562226 345774 562294
rect 345154 562170 345250 562226
rect 345306 562170 345374 562226
rect 345430 562170 345498 562226
rect 345554 562170 345622 562226
rect 345678 562170 345774 562226
rect 345154 562102 345774 562170
rect 345154 562046 345250 562102
rect 345306 562046 345374 562102
rect 345430 562046 345498 562102
rect 345554 562046 345622 562102
rect 345678 562046 345774 562102
rect 345154 561978 345774 562046
rect 345154 561922 345250 561978
rect 345306 561922 345374 561978
rect 345430 561922 345498 561978
rect 345554 561922 345622 561978
rect 345678 561922 345774 561978
rect 345154 544350 345774 561922
rect 345154 544294 345250 544350
rect 345306 544294 345374 544350
rect 345430 544294 345498 544350
rect 345554 544294 345622 544350
rect 345678 544294 345774 544350
rect 345154 544226 345774 544294
rect 345154 544170 345250 544226
rect 345306 544170 345374 544226
rect 345430 544170 345498 544226
rect 345554 544170 345622 544226
rect 345678 544170 345774 544226
rect 345154 544102 345774 544170
rect 345154 544046 345250 544102
rect 345306 544046 345374 544102
rect 345430 544046 345498 544102
rect 345554 544046 345622 544102
rect 345678 544046 345774 544102
rect 345154 543978 345774 544046
rect 345154 543922 345250 543978
rect 345306 543922 345374 543978
rect 345430 543922 345498 543978
rect 345554 543922 345622 543978
rect 345678 543922 345774 543978
rect 345154 527750 345774 543922
rect 348874 598172 349494 598268
rect 348874 598116 348970 598172
rect 349026 598116 349094 598172
rect 349150 598116 349218 598172
rect 349274 598116 349342 598172
rect 349398 598116 349494 598172
rect 348874 598048 349494 598116
rect 348874 597992 348970 598048
rect 349026 597992 349094 598048
rect 349150 597992 349218 598048
rect 349274 597992 349342 598048
rect 349398 597992 349494 598048
rect 348874 597924 349494 597992
rect 348874 597868 348970 597924
rect 349026 597868 349094 597924
rect 349150 597868 349218 597924
rect 349274 597868 349342 597924
rect 349398 597868 349494 597924
rect 348874 597800 349494 597868
rect 348874 597744 348970 597800
rect 349026 597744 349094 597800
rect 349150 597744 349218 597800
rect 349274 597744 349342 597800
rect 349398 597744 349494 597800
rect 348874 586350 349494 597744
rect 348874 586294 348970 586350
rect 349026 586294 349094 586350
rect 349150 586294 349218 586350
rect 349274 586294 349342 586350
rect 349398 586294 349494 586350
rect 348874 586226 349494 586294
rect 348874 586170 348970 586226
rect 349026 586170 349094 586226
rect 349150 586170 349218 586226
rect 349274 586170 349342 586226
rect 349398 586170 349494 586226
rect 348874 586102 349494 586170
rect 348874 586046 348970 586102
rect 349026 586046 349094 586102
rect 349150 586046 349218 586102
rect 349274 586046 349342 586102
rect 349398 586046 349494 586102
rect 348874 585978 349494 586046
rect 348874 585922 348970 585978
rect 349026 585922 349094 585978
rect 349150 585922 349218 585978
rect 349274 585922 349342 585978
rect 349398 585922 349494 585978
rect 348874 568350 349494 585922
rect 348874 568294 348970 568350
rect 349026 568294 349094 568350
rect 349150 568294 349218 568350
rect 349274 568294 349342 568350
rect 349398 568294 349494 568350
rect 348874 568226 349494 568294
rect 348874 568170 348970 568226
rect 349026 568170 349094 568226
rect 349150 568170 349218 568226
rect 349274 568170 349342 568226
rect 349398 568170 349494 568226
rect 348874 568102 349494 568170
rect 348874 568046 348970 568102
rect 349026 568046 349094 568102
rect 349150 568046 349218 568102
rect 349274 568046 349342 568102
rect 349398 568046 349494 568102
rect 348874 567978 349494 568046
rect 348874 567922 348970 567978
rect 349026 567922 349094 567978
rect 349150 567922 349218 567978
rect 349274 567922 349342 567978
rect 349398 567922 349494 567978
rect 348874 550350 349494 567922
rect 348874 550294 348970 550350
rect 349026 550294 349094 550350
rect 349150 550294 349218 550350
rect 349274 550294 349342 550350
rect 349398 550294 349494 550350
rect 348874 550226 349494 550294
rect 348874 550170 348970 550226
rect 349026 550170 349094 550226
rect 349150 550170 349218 550226
rect 349274 550170 349342 550226
rect 349398 550170 349494 550226
rect 348874 550102 349494 550170
rect 348874 550046 348970 550102
rect 349026 550046 349094 550102
rect 349150 550046 349218 550102
rect 349274 550046 349342 550102
rect 349398 550046 349494 550102
rect 348874 549978 349494 550046
rect 348874 549922 348970 549978
rect 349026 549922 349094 549978
rect 349150 549922 349218 549978
rect 349274 549922 349342 549978
rect 349398 549922 349494 549978
rect 348874 532350 349494 549922
rect 348874 532294 348970 532350
rect 349026 532294 349094 532350
rect 349150 532294 349218 532350
rect 349274 532294 349342 532350
rect 349398 532294 349494 532350
rect 348874 532226 349494 532294
rect 348874 532170 348970 532226
rect 349026 532170 349094 532226
rect 349150 532170 349218 532226
rect 349274 532170 349342 532226
rect 349398 532170 349494 532226
rect 348874 532102 349494 532170
rect 348874 532046 348970 532102
rect 349026 532046 349094 532102
rect 349150 532046 349218 532102
rect 349274 532046 349342 532102
rect 349398 532046 349494 532102
rect 348874 531978 349494 532046
rect 348874 531922 348970 531978
rect 349026 531922 349094 531978
rect 349150 531922 349218 531978
rect 349274 531922 349342 531978
rect 349398 531922 349494 531978
rect 348874 527750 349494 531922
rect 363154 597212 363774 598268
rect 363154 597156 363250 597212
rect 363306 597156 363374 597212
rect 363430 597156 363498 597212
rect 363554 597156 363622 597212
rect 363678 597156 363774 597212
rect 363154 597088 363774 597156
rect 363154 597032 363250 597088
rect 363306 597032 363374 597088
rect 363430 597032 363498 597088
rect 363554 597032 363622 597088
rect 363678 597032 363774 597088
rect 363154 596964 363774 597032
rect 363154 596908 363250 596964
rect 363306 596908 363374 596964
rect 363430 596908 363498 596964
rect 363554 596908 363622 596964
rect 363678 596908 363774 596964
rect 363154 596840 363774 596908
rect 363154 596784 363250 596840
rect 363306 596784 363374 596840
rect 363430 596784 363498 596840
rect 363554 596784 363622 596840
rect 363678 596784 363774 596840
rect 363154 580350 363774 596784
rect 363154 580294 363250 580350
rect 363306 580294 363374 580350
rect 363430 580294 363498 580350
rect 363554 580294 363622 580350
rect 363678 580294 363774 580350
rect 363154 580226 363774 580294
rect 363154 580170 363250 580226
rect 363306 580170 363374 580226
rect 363430 580170 363498 580226
rect 363554 580170 363622 580226
rect 363678 580170 363774 580226
rect 363154 580102 363774 580170
rect 363154 580046 363250 580102
rect 363306 580046 363374 580102
rect 363430 580046 363498 580102
rect 363554 580046 363622 580102
rect 363678 580046 363774 580102
rect 363154 579978 363774 580046
rect 363154 579922 363250 579978
rect 363306 579922 363374 579978
rect 363430 579922 363498 579978
rect 363554 579922 363622 579978
rect 363678 579922 363774 579978
rect 363154 562350 363774 579922
rect 363154 562294 363250 562350
rect 363306 562294 363374 562350
rect 363430 562294 363498 562350
rect 363554 562294 363622 562350
rect 363678 562294 363774 562350
rect 363154 562226 363774 562294
rect 363154 562170 363250 562226
rect 363306 562170 363374 562226
rect 363430 562170 363498 562226
rect 363554 562170 363622 562226
rect 363678 562170 363774 562226
rect 363154 562102 363774 562170
rect 363154 562046 363250 562102
rect 363306 562046 363374 562102
rect 363430 562046 363498 562102
rect 363554 562046 363622 562102
rect 363678 562046 363774 562102
rect 363154 561978 363774 562046
rect 363154 561922 363250 561978
rect 363306 561922 363374 561978
rect 363430 561922 363498 561978
rect 363554 561922 363622 561978
rect 363678 561922 363774 561978
rect 363154 544350 363774 561922
rect 363154 544294 363250 544350
rect 363306 544294 363374 544350
rect 363430 544294 363498 544350
rect 363554 544294 363622 544350
rect 363678 544294 363774 544350
rect 363154 544226 363774 544294
rect 363154 544170 363250 544226
rect 363306 544170 363374 544226
rect 363430 544170 363498 544226
rect 363554 544170 363622 544226
rect 363678 544170 363774 544226
rect 363154 544102 363774 544170
rect 363154 544046 363250 544102
rect 363306 544046 363374 544102
rect 363430 544046 363498 544102
rect 363554 544046 363622 544102
rect 363678 544046 363774 544102
rect 363154 543978 363774 544046
rect 363154 543922 363250 543978
rect 363306 543922 363374 543978
rect 363430 543922 363498 543978
rect 363554 543922 363622 543978
rect 363678 543922 363774 543978
rect 363154 527750 363774 543922
rect 366874 598172 367494 598268
rect 366874 598116 366970 598172
rect 367026 598116 367094 598172
rect 367150 598116 367218 598172
rect 367274 598116 367342 598172
rect 367398 598116 367494 598172
rect 366874 598048 367494 598116
rect 366874 597992 366970 598048
rect 367026 597992 367094 598048
rect 367150 597992 367218 598048
rect 367274 597992 367342 598048
rect 367398 597992 367494 598048
rect 366874 597924 367494 597992
rect 366874 597868 366970 597924
rect 367026 597868 367094 597924
rect 367150 597868 367218 597924
rect 367274 597868 367342 597924
rect 367398 597868 367494 597924
rect 366874 597800 367494 597868
rect 366874 597744 366970 597800
rect 367026 597744 367094 597800
rect 367150 597744 367218 597800
rect 367274 597744 367342 597800
rect 367398 597744 367494 597800
rect 366874 586350 367494 597744
rect 366874 586294 366970 586350
rect 367026 586294 367094 586350
rect 367150 586294 367218 586350
rect 367274 586294 367342 586350
rect 367398 586294 367494 586350
rect 366874 586226 367494 586294
rect 366874 586170 366970 586226
rect 367026 586170 367094 586226
rect 367150 586170 367218 586226
rect 367274 586170 367342 586226
rect 367398 586170 367494 586226
rect 366874 586102 367494 586170
rect 366874 586046 366970 586102
rect 367026 586046 367094 586102
rect 367150 586046 367218 586102
rect 367274 586046 367342 586102
rect 367398 586046 367494 586102
rect 366874 585978 367494 586046
rect 366874 585922 366970 585978
rect 367026 585922 367094 585978
rect 367150 585922 367218 585978
rect 367274 585922 367342 585978
rect 367398 585922 367494 585978
rect 366874 568350 367494 585922
rect 366874 568294 366970 568350
rect 367026 568294 367094 568350
rect 367150 568294 367218 568350
rect 367274 568294 367342 568350
rect 367398 568294 367494 568350
rect 366874 568226 367494 568294
rect 366874 568170 366970 568226
rect 367026 568170 367094 568226
rect 367150 568170 367218 568226
rect 367274 568170 367342 568226
rect 367398 568170 367494 568226
rect 366874 568102 367494 568170
rect 366874 568046 366970 568102
rect 367026 568046 367094 568102
rect 367150 568046 367218 568102
rect 367274 568046 367342 568102
rect 367398 568046 367494 568102
rect 366874 567978 367494 568046
rect 366874 567922 366970 567978
rect 367026 567922 367094 567978
rect 367150 567922 367218 567978
rect 367274 567922 367342 567978
rect 367398 567922 367494 567978
rect 366874 550350 367494 567922
rect 366874 550294 366970 550350
rect 367026 550294 367094 550350
rect 367150 550294 367218 550350
rect 367274 550294 367342 550350
rect 367398 550294 367494 550350
rect 366874 550226 367494 550294
rect 366874 550170 366970 550226
rect 367026 550170 367094 550226
rect 367150 550170 367218 550226
rect 367274 550170 367342 550226
rect 367398 550170 367494 550226
rect 366874 550102 367494 550170
rect 366874 550046 366970 550102
rect 367026 550046 367094 550102
rect 367150 550046 367218 550102
rect 367274 550046 367342 550102
rect 367398 550046 367494 550102
rect 366874 549978 367494 550046
rect 366874 549922 366970 549978
rect 367026 549922 367094 549978
rect 367150 549922 367218 549978
rect 367274 549922 367342 549978
rect 367398 549922 367494 549978
rect 366874 532350 367494 549922
rect 366874 532294 366970 532350
rect 367026 532294 367094 532350
rect 367150 532294 367218 532350
rect 367274 532294 367342 532350
rect 367398 532294 367494 532350
rect 366874 532226 367494 532294
rect 366874 532170 366970 532226
rect 367026 532170 367094 532226
rect 367150 532170 367218 532226
rect 367274 532170 367342 532226
rect 367398 532170 367494 532226
rect 366874 532102 367494 532170
rect 366874 532046 366970 532102
rect 367026 532046 367094 532102
rect 367150 532046 367218 532102
rect 367274 532046 367342 532102
rect 367398 532046 367494 532102
rect 366874 531978 367494 532046
rect 366874 531922 366970 531978
rect 367026 531922 367094 531978
rect 367150 531922 367218 531978
rect 367274 531922 367342 531978
rect 367398 531922 367494 531978
rect 366874 527750 367494 531922
rect 381154 597212 381774 598268
rect 381154 597156 381250 597212
rect 381306 597156 381374 597212
rect 381430 597156 381498 597212
rect 381554 597156 381622 597212
rect 381678 597156 381774 597212
rect 381154 597088 381774 597156
rect 381154 597032 381250 597088
rect 381306 597032 381374 597088
rect 381430 597032 381498 597088
rect 381554 597032 381622 597088
rect 381678 597032 381774 597088
rect 381154 596964 381774 597032
rect 381154 596908 381250 596964
rect 381306 596908 381374 596964
rect 381430 596908 381498 596964
rect 381554 596908 381622 596964
rect 381678 596908 381774 596964
rect 381154 596840 381774 596908
rect 381154 596784 381250 596840
rect 381306 596784 381374 596840
rect 381430 596784 381498 596840
rect 381554 596784 381622 596840
rect 381678 596784 381774 596840
rect 381154 580350 381774 596784
rect 381154 580294 381250 580350
rect 381306 580294 381374 580350
rect 381430 580294 381498 580350
rect 381554 580294 381622 580350
rect 381678 580294 381774 580350
rect 381154 580226 381774 580294
rect 381154 580170 381250 580226
rect 381306 580170 381374 580226
rect 381430 580170 381498 580226
rect 381554 580170 381622 580226
rect 381678 580170 381774 580226
rect 381154 580102 381774 580170
rect 381154 580046 381250 580102
rect 381306 580046 381374 580102
rect 381430 580046 381498 580102
rect 381554 580046 381622 580102
rect 381678 580046 381774 580102
rect 381154 579978 381774 580046
rect 381154 579922 381250 579978
rect 381306 579922 381374 579978
rect 381430 579922 381498 579978
rect 381554 579922 381622 579978
rect 381678 579922 381774 579978
rect 381154 562350 381774 579922
rect 381154 562294 381250 562350
rect 381306 562294 381374 562350
rect 381430 562294 381498 562350
rect 381554 562294 381622 562350
rect 381678 562294 381774 562350
rect 381154 562226 381774 562294
rect 381154 562170 381250 562226
rect 381306 562170 381374 562226
rect 381430 562170 381498 562226
rect 381554 562170 381622 562226
rect 381678 562170 381774 562226
rect 381154 562102 381774 562170
rect 381154 562046 381250 562102
rect 381306 562046 381374 562102
rect 381430 562046 381498 562102
rect 381554 562046 381622 562102
rect 381678 562046 381774 562102
rect 381154 561978 381774 562046
rect 381154 561922 381250 561978
rect 381306 561922 381374 561978
rect 381430 561922 381498 561978
rect 381554 561922 381622 561978
rect 381678 561922 381774 561978
rect 381154 544350 381774 561922
rect 381154 544294 381250 544350
rect 381306 544294 381374 544350
rect 381430 544294 381498 544350
rect 381554 544294 381622 544350
rect 381678 544294 381774 544350
rect 381154 544226 381774 544294
rect 381154 544170 381250 544226
rect 381306 544170 381374 544226
rect 381430 544170 381498 544226
rect 381554 544170 381622 544226
rect 381678 544170 381774 544226
rect 381154 544102 381774 544170
rect 381154 544046 381250 544102
rect 381306 544046 381374 544102
rect 381430 544046 381498 544102
rect 381554 544046 381622 544102
rect 381678 544046 381774 544102
rect 381154 543978 381774 544046
rect 381154 543922 381250 543978
rect 381306 543922 381374 543978
rect 381430 543922 381498 543978
rect 381554 543922 381622 543978
rect 381678 543922 381774 543978
rect 381154 527750 381774 543922
rect 384874 598172 385494 598268
rect 384874 598116 384970 598172
rect 385026 598116 385094 598172
rect 385150 598116 385218 598172
rect 385274 598116 385342 598172
rect 385398 598116 385494 598172
rect 384874 598048 385494 598116
rect 384874 597992 384970 598048
rect 385026 597992 385094 598048
rect 385150 597992 385218 598048
rect 385274 597992 385342 598048
rect 385398 597992 385494 598048
rect 384874 597924 385494 597992
rect 384874 597868 384970 597924
rect 385026 597868 385094 597924
rect 385150 597868 385218 597924
rect 385274 597868 385342 597924
rect 385398 597868 385494 597924
rect 384874 597800 385494 597868
rect 384874 597744 384970 597800
rect 385026 597744 385094 597800
rect 385150 597744 385218 597800
rect 385274 597744 385342 597800
rect 385398 597744 385494 597800
rect 384874 586350 385494 597744
rect 384874 586294 384970 586350
rect 385026 586294 385094 586350
rect 385150 586294 385218 586350
rect 385274 586294 385342 586350
rect 385398 586294 385494 586350
rect 384874 586226 385494 586294
rect 384874 586170 384970 586226
rect 385026 586170 385094 586226
rect 385150 586170 385218 586226
rect 385274 586170 385342 586226
rect 385398 586170 385494 586226
rect 384874 586102 385494 586170
rect 384874 586046 384970 586102
rect 385026 586046 385094 586102
rect 385150 586046 385218 586102
rect 385274 586046 385342 586102
rect 385398 586046 385494 586102
rect 384874 585978 385494 586046
rect 384874 585922 384970 585978
rect 385026 585922 385094 585978
rect 385150 585922 385218 585978
rect 385274 585922 385342 585978
rect 385398 585922 385494 585978
rect 384874 568350 385494 585922
rect 384874 568294 384970 568350
rect 385026 568294 385094 568350
rect 385150 568294 385218 568350
rect 385274 568294 385342 568350
rect 385398 568294 385494 568350
rect 384874 568226 385494 568294
rect 384874 568170 384970 568226
rect 385026 568170 385094 568226
rect 385150 568170 385218 568226
rect 385274 568170 385342 568226
rect 385398 568170 385494 568226
rect 384874 568102 385494 568170
rect 384874 568046 384970 568102
rect 385026 568046 385094 568102
rect 385150 568046 385218 568102
rect 385274 568046 385342 568102
rect 385398 568046 385494 568102
rect 384874 567978 385494 568046
rect 384874 567922 384970 567978
rect 385026 567922 385094 567978
rect 385150 567922 385218 567978
rect 385274 567922 385342 567978
rect 385398 567922 385494 567978
rect 384874 550350 385494 567922
rect 384874 550294 384970 550350
rect 385026 550294 385094 550350
rect 385150 550294 385218 550350
rect 385274 550294 385342 550350
rect 385398 550294 385494 550350
rect 384874 550226 385494 550294
rect 384874 550170 384970 550226
rect 385026 550170 385094 550226
rect 385150 550170 385218 550226
rect 385274 550170 385342 550226
rect 385398 550170 385494 550226
rect 384874 550102 385494 550170
rect 384874 550046 384970 550102
rect 385026 550046 385094 550102
rect 385150 550046 385218 550102
rect 385274 550046 385342 550102
rect 385398 550046 385494 550102
rect 384874 549978 385494 550046
rect 384874 549922 384970 549978
rect 385026 549922 385094 549978
rect 385150 549922 385218 549978
rect 385274 549922 385342 549978
rect 385398 549922 385494 549978
rect 384874 532350 385494 549922
rect 384874 532294 384970 532350
rect 385026 532294 385094 532350
rect 385150 532294 385218 532350
rect 385274 532294 385342 532350
rect 385398 532294 385494 532350
rect 384874 532226 385494 532294
rect 384874 532170 384970 532226
rect 385026 532170 385094 532226
rect 385150 532170 385218 532226
rect 385274 532170 385342 532226
rect 385398 532170 385494 532226
rect 384874 532102 385494 532170
rect 384874 532046 384970 532102
rect 385026 532046 385094 532102
rect 385150 532046 385218 532102
rect 385274 532046 385342 532102
rect 385398 532046 385494 532102
rect 384874 531978 385494 532046
rect 384874 531922 384970 531978
rect 385026 531922 385094 531978
rect 385150 531922 385218 531978
rect 385274 531922 385342 531978
rect 385398 531922 385494 531978
rect 384874 527750 385494 531922
rect 399154 597212 399774 598268
rect 399154 597156 399250 597212
rect 399306 597156 399374 597212
rect 399430 597156 399498 597212
rect 399554 597156 399622 597212
rect 399678 597156 399774 597212
rect 399154 597088 399774 597156
rect 399154 597032 399250 597088
rect 399306 597032 399374 597088
rect 399430 597032 399498 597088
rect 399554 597032 399622 597088
rect 399678 597032 399774 597088
rect 399154 596964 399774 597032
rect 399154 596908 399250 596964
rect 399306 596908 399374 596964
rect 399430 596908 399498 596964
rect 399554 596908 399622 596964
rect 399678 596908 399774 596964
rect 399154 596840 399774 596908
rect 399154 596784 399250 596840
rect 399306 596784 399374 596840
rect 399430 596784 399498 596840
rect 399554 596784 399622 596840
rect 399678 596784 399774 596840
rect 399154 580350 399774 596784
rect 399154 580294 399250 580350
rect 399306 580294 399374 580350
rect 399430 580294 399498 580350
rect 399554 580294 399622 580350
rect 399678 580294 399774 580350
rect 399154 580226 399774 580294
rect 399154 580170 399250 580226
rect 399306 580170 399374 580226
rect 399430 580170 399498 580226
rect 399554 580170 399622 580226
rect 399678 580170 399774 580226
rect 399154 580102 399774 580170
rect 399154 580046 399250 580102
rect 399306 580046 399374 580102
rect 399430 580046 399498 580102
rect 399554 580046 399622 580102
rect 399678 580046 399774 580102
rect 399154 579978 399774 580046
rect 399154 579922 399250 579978
rect 399306 579922 399374 579978
rect 399430 579922 399498 579978
rect 399554 579922 399622 579978
rect 399678 579922 399774 579978
rect 399154 562350 399774 579922
rect 399154 562294 399250 562350
rect 399306 562294 399374 562350
rect 399430 562294 399498 562350
rect 399554 562294 399622 562350
rect 399678 562294 399774 562350
rect 399154 562226 399774 562294
rect 399154 562170 399250 562226
rect 399306 562170 399374 562226
rect 399430 562170 399498 562226
rect 399554 562170 399622 562226
rect 399678 562170 399774 562226
rect 399154 562102 399774 562170
rect 399154 562046 399250 562102
rect 399306 562046 399374 562102
rect 399430 562046 399498 562102
rect 399554 562046 399622 562102
rect 399678 562046 399774 562102
rect 399154 561978 399774 562046
rect 399154 561922 399250 561978
rect 399306 561922 399374 561978
rect 399430 561922 399498 561978
rect 399554 561922 399622 561978
rect 399678 561922 399774 561978
rect 399154 544350 399774 561922
rect 399154 544294 399250 544350
rect 399306 544294 399374 544350
rect 399430 544294 399498 544350
rect 399554 544294 399622 544350
rect 399678 544294 399774 544350
rect 399154 544226 399774 544294
rect 399154 544170 399250 544226
rect 399306 544170 399374 544226
rect 399430 544170 399498 544226
rect 399554 544170 399622 544226
rect 399678 544170 399774 544226
rect 399154 544102 399774 544170
rect 399154 544046 399250 544102
rect 399306 544046 399374 544102
rect 399430 544046 399498 544102
rect 399554 544046 399622 544102
rect 399678 544046 399774 544102
rect 399154 543978 399774 544046
rect 399154 543922 399250 543978
rect 399306 543922 399374 543978
rect 399430 543922 399498 543978
rect 399554 543922 399622 543978
rect 399678 543922 399774 543978
rect 399154 527750 399774 543922
rect 402874 598172 403494 598268
rect 402874 598116 402970 598172
rect 403026 598116 403094 598172
rect 403150 598116 403218 598172
rect 403274 598116 403342 598172
rect 403398 598116 403494 598172
rect 402874 598048 403494 598116
rect 402874 597992 402970 598048
rect 403026 597992 403094 598048
rect 403150 597992 403218 598048
rect 403274 597992 403342 598048
rect 403398 597992 403494 598048
rect 402874 597924 403494 597992
rect 402874 597868 402970 597924
rect 403026 597868 403094 597924
rect 403150 597868 403218 597924
rect 403274 597868 403342 597924
rect 403398 597868 403494 597924
rect 402874 597800 403494 597868
rect 402874 597744 402970 597800
rect 403026 597744 403094 597800
rect 403150 597744 403218 597800
rect 403274 597744 403342 597800
rect 403398 597744 403494 597800
rect 402874 586350 403494 597744
rect 402874 586294 402970 586350
rect 403026 586294 403094 586350
rect 403150 586294 403218 586350
rect 403274 586294 403342 586350
rect 403398 586294 403494 586350
rect 402874 586226 403494 586294
rect 402874 586170 402970 586226
rect 403026 586170 403094 586226
rect 403150 586170 403218 586226
rect 403274 586170 403342 586226
rect 403398 586170 403494 586226
rect 402874 586102 403494 586170
rect 402874 586046 402970 586102
rect 403026 586046 403094 586102
rect 403150 586046 403218 586102
rect 403274 586046 403342 586102
rect 403398 586046 403494 586102
rect 402874 585978 403494 586046
rect 402874 585922 402970 585978
rect 403026 585922 403094 585978
rect 403150 585922 403218 585978
rect 403274 585922 403342 585978
rect 403398 585922 403494 585978
rect 402874 568350 403494 585922
rect 402874 568294 402970 568350
rect 403026 568294 403094 568350
rect 403150 568294 403218 568350
rect 403274 568294 403342 568350
rect 403398 568294 403494 568350
rect 402874 568226 403494 568294
rect 402874 568170 402970 568226
rect 403026 568170 403094 568226
rect 403150 568170 403218 568226
rect 403274 568170 403342 568226
rect 403398 568170 403494 568226
rect 402874 568102 403494 568170
rect 402874 568046 402970 568102
rect 403026 568046 403094 568102
rect 403150 568046 403218 568102
rect 403274 568046 403342 568102
rect 403398 568046 403494 568102
rect 402874 567978 403494 568046
rect 402874 567922 402970 567978
rect 403026 567922 403094 567978
rect 403150 567922 403218 567978
rect 403274 567922 403342 567978
rect 403398 567922 403494 567978
rect 402874 550350 403494 567922
rect 402874 550294 402970 550350
rect 403026 550294 403094 550350
rect 403150 550294 403218 550350
rect 403274 550294 403342 550350
rect 403398 550294 403494 550350
rect 402874 550226 403494 550294
rect 402874 550170 402970 550226
rect 403026 550170 403094 550226
rect 403150 550170 403218 550226
rect 403274 550170 403342 550226
rect 403398 550170 403494 550226
rect 402874 550102 403494 550170
rect 402874 550046 402970 550102
rect 403026 550046 403094 550102
rect 403150 550046 403218 550102
rect 403274 550046 403342 550102
rect 403398 550046 403494 550102
rect 402874 549978 403494 550046
rect 402874 549922 402970 549978
rect 403026 549922 403094 549978
rect 403150 549922 403218 549978
rect 403274 549922 403342 549978
rect 403398 549922 403494 549978
rect 402874 532350 403494 549922
rect 402874 532294 402970 532350
rect 403026 532294 403094 532350
rect 403150 532294 403218 532350
rect 403274 532294 403342 532350
rect 403398 532294 403494 532350
rect 402874 532226 403494 532294
rect 402874 532170 402970 532226
rect 403026 532170 403094 532226
rect 403150 532170 403218 532226
rect 403274 532170 403342 532226
rect 403398 532170 403494 532226
rect 402874 532102 403494 532170
rect 402874 532046 402970 532102
rect 403026 532046 403094 532102
rect 403150 532046 403218 532102
rect 403274 532046 403342 532102
rect 403398 532046 403494 532102
rect 402874 531978 403494 532046
rect 402874 531922 402970 531978
rect 403026 531922 403094 531978
rect 403150 531922 403218 531978
rect 403274 531922 403342 531978
rect 403398 531922 403494 531978
rect 402874 527750 403494 531922
rect 417154 597212 417774 598268
rect 417154 597156 417250 597212
rect 417306 597156 417374 597212
rect 417430 597156 417498 597212
rect 417554 597156 417622 597212
rect 417678 597156 417774 597212
rect 417154 597088 417774 597156
rect 417154 597032 417250 597088
rect 417306 597032 417374 597088
rect 417430 597032 417498 597088
rect 417554 597032 417622 597088
rect 417678 597032 417774 597088
rect 417154 596964 417774 597032
rect 417154 596908 417250 596964
rect 417306 596908 417374 596964
rect 417430 596908 417498 596964
rect 417554 596908 417622 596964
rect 417678 596908 417774 596964
rect 417154 596840 417774 596908
rect 417154 596784 417250 596840
rect 417306 596784 417374 596840
rect 417430 596784 417498 596840
rect 417554 596784 417622 596840
rect 417678 596784 417774 596840
rect 417154 580350 417774 596784
rect 417154 580294 417250 580350
rect 417306 580294 417374 580350
rect 417430 580294 417498 580350
rect 417554 580294 417622 580350
rect 417678 580294 417774 580350
rect 417154 580226 417774 580294
rect 417154 580170 417250 580226
rect 417306 580170 417374 580226
rect 417430 580170 417498 580226
rect 417554 580170 417622 580226
rect 417678 580170 417774 580226
rect 417154 580102 417774 580170
rect 417154 580046 417250 580102
rect 417306 580046 417374 580102
rect 417430 580046 417498 580102
rect 417554 580046 417622 580102
rect 417678 580046 417774 580102
rect 417154 579978 417774 580046
rect 417154 579922 417250 579978
rect 417306 579922 417374 579978
rect 417430 579922 417498 579978
rect 417554 579922 417622 579978
rect 417678 579922 417774 579978
rect 417154 562350 417774 579922
rect 417154 562294 417250 562350
rect 417306 562294 417374 562350
rect 417430 562294 417498 562350
rect 417554 562294 417622 562350
rect 417678 562294 417774 562350
rect 417154 562226 417774 562294
rect 417154 562170 417250 562226
rect 417306 562170 417374 562226
rect 417430 562170 417498 562226
rect 417554 562170 417622 562226
rect 417678 562170 417774 562226
rect 417154 562102 417774 562170
rect 417154 562046 417250 562102
rect 417306 562046 417374 562102
rect 417430 562046 417498 562102
rect 417554 562046 417622 562102
rect 417678 562046 417774 562102
rect 417154 561978 417774 562046
rect 417154 561922 417250 561978
rect 417306 561922 417374 561978
rect 417430 561922 417498 561978
rect 417554 561922 417622 561978
rect 417678 561922 417774 561978
rect 417154 544350 417774 561922
rect 417154 544294 417250 544350
rect 417306 544294 417374 544350
rect 417430 544294 417498 544350
rect 417554 544294 417622 544350
rect 417678 544294 417774 544350
rect 417154 544226 417774 544294
rect 417154 544170 417250 544226
rect 417306 544170 417374 544226
rect 417430 544170 417498 544226
rect 417554 544170 417622 544226
rect 417678 544170 417774 544226
rect 417154 544102 417774 544170
rect 417154 544046 417250 544102
rect 417306 544046 417374 544102
rect 417430 544046 417498 544102
rect 417554 544046 417622 544102
rect 417678 544046 417774 544102
rect 417154 543978 417774 544046
rect 417154 543922 417250 543978
rect 417306 543922 417374 543978
rect 417430 543922 417498 543978
rect 417554 543922 417622 543978
rect 417678 543922 417774 543978
rect 417154 527750 417774 543922
rect 420874 598172 421494 598268
rect 420874 598116 420970 598172
rect 421026 598116 421094 598172
rect 421150 598116 421218 598172
rect 421274 598116 421342 598172
rect 421398 598116 421494 598172
rect 420874 598048 421494 598116
rect 420874 597992 420970 598048
rect 421026 597992 421094 598048
rect 421150 597992 421218 598048
rect 421274 597992 421342 598048
rect 421398 597992 421494 598048
rect 420874 597924 421494 597992
rect 420874 597868 420970 597924
rect 421026 597868 421094 597924
rect 421150 597868 421218 597924
rect 421274 597868 421342 597924
rect 421398 597868 421494 597924
rect 420874 597800 421494 597868
rect 420874 597744 420970 597800
rect 421026 597744 421094 597800
rect 421150 597744 421218 597800
rect 421274 597744 421342 597800
rect 421398 597744 421494 597800
rect 420874 586350 421494 597744
rect 420874 586294 420970 586350
rect 421026 586294 421094 586350
rect 421150 586294 421218 586350
rect 421274 586294 421342 586350
rect 421398 586294 421494 586350
rect 420874 586226 421494 586294
rect 420874 586170 420970 586226
rect 421026 586170 421094 586226
rect 421150 586170 421218 586226
rect 421274 586170 421342 586226
rect 421398 586170 421494 586226
rect 420874 586102 421494 586170
rect 420874 586046 420970 586102
rect 421026 586046 421094 586102
rect 421150 586046 421218 586102
rect 421274 586046 421342 586102
rect 421398 586046 421494 586102
rect 420874 585978 421494 586046
rect 420874 585922 420970 585978
rect 421026 585922 421094 585978
rect 421150 585922 421218 585978
rect 421274 585922 421342 585978
rect 421398 585922 421494 585978
rect 420874 568350 421494 585922
rect 420874 568294 420970 568350
rect 421026 568294 421094 568350
rect 421150 568294 421218 568350
rect 421274 568294 421342 568350
rect 421398 568294 421494 568350
rect 420874 568226 421494 568294
rect 420874 568170 420970 568226
rect 421026 568170 421094 568226
rect 421150 568170 421218 568226
rect 421274 568170 421342 568226
rect 421398 568170 421494 568226
rect 420874 568102 421494 568170
rect 420874 568046 420970 568102
rect 421026 568046 421094 568102
rect 421150 568046 421218 568102
rect 421274 568046 421342 568102
rect 421398 568046 421494 568102
rect 420874 567978 421494 568046
rect 420874 567922 420970 567978
rect 421026 567922 421094 567978
rect 421150 567922 421218 567978
rect 421274 567922 421342 567978
rect 421398 567922 421494 567978
rect 420874 550350 421494 567922
rect 420874 550294 420970 550350
rect 421026 550294 421094 550350
rect 421150 550294 421218 550350
rect 421274 550294 421342 550350
rect 421398 550294 421494 550350
rect 420874 550226 421494 550294
rect 420874 550170 420970 550226
rect 421026 550170 421094 550226
rect 421150 550170 421218 550226
rect 421274 550170 421342 550226
rect 421398 550170 421494 550226
rect 420874 550102 421494 550170
rect 420874 550046 420970 550102
rect 421026 550046 421094 550102
rect 421150 550046 421218 550102
rect 421274 550046 421342 550102
rect 421398 550046 421494 550102
rect 420874 549978 421494 550046
rect 420874 549922 420970 549978
rect 421026 549922 421094 549978
rect 421150 549922 421218 549978
rect 421274 549922 421342 549978
rect 421398 549922 421494 549978
rect 420874 532350 421494 549922
rect 420874 532294 420970 532350
rect 421026 532294 421094 532350
rect 421150 532294 421218 532350
rect 421274 532294 421342 532350
rect 421398 532294 421494 532350
rect 420874 532226 421494 532294
rect 420874 532170 420970 532226
rect 421026 532170 421094 532226
rect 421150 532170 421218 532226
rect 421274 532170 421342 532226
rect 421398 532170 421494 532226
rect 420874 532102 421494 532170
rect 420874 532046 420970 532102
rect 421026 532046 421094 532102
rect 421150 532046 421218 532102
rect 421274 532046 421342 532102
rect 421398 532046 421494 532102
rect 420874 531978 421494 532046
rect 420874 531922 420970 531978
rect 421026 531922 421094 531978
rect 421150 531922 421218 531978
rect 421274 531922 421342 531978
rect 421398 531922 421494 531978
rect 420874 527750 421494 531922
rect 435154 597212 435774 598268
rect 435154 597156 435250 597212
rect 435306 597156 435374 597212
rect 435430 597156 435498 597212
rect 435554 597156 435622 597212
rect 435678 597156 435774 597212
rect 435154 597088 435774 597156
rect 435154 597032 435250 597088
rect 435306 597032 435374 597088
rect 435430 597032 435498 597088
rect 435554 597032 435622 597088
rect 435678 597032 435774 597088
rect 435154 596964 435774 597032
rect 435154 596908 435250 596964
rect 435306 596908 435374 596964
rect 435430 596908 435498 596964
rect 435554 596908 435622 596964
rect 435678 596908 435774 596964
rect 435154 596840 435774 596908
rect 435154 596784 435250 596840
rect 435306 596784 435374 596840
rect 435430 596784 435498 596840
rect 435554 596784 435622 596840
rect 435678 596784 435774 596840
rect 435154 580350 435774 596784
rect 435154 580294 435250 580350
rect 435306 580294 435374 580350
rect 435430 580294 435498 580350
rect 435554 580294 435622 580350
rect 435678 580294 435774 580350
rect 435154 580226 435774 580294
rect 435154 580170 435250 580226
rect 435306 580170 435374 580226
rect 435430 580170 435498 580226
rect 435554 580170 435622 580226
rect 435678 580170 435774 580226
rect 435154 580102 435774 580170
rect 435154 580046 435250 580102
rect 435306 580046 435374 580102
rect 435430 580046 435498 580102
rect 435554 580046 435622 580102
rect 435678 580046 435774 580102
rect 435154 579978 435774 580046
rect 435154 579922 435250 579978
rect 435306 579922 435374 579978
rect 435430 579922 435498 579978
rect 435554 579922 435622 579978
rect 435678 579922 435774 579978
rect 435154 562350 435774 579922
rect 435154 562294 435250 562350
rect 435306 562294 435374 562350
rect 435430 562294 435498 562350
rect 435554 562294 435622 562350
rect 435678 562294 435774 562350
rect 435154 562226 435774 562294
rect 435154 562170 435250 562226
rect 435306 562170 435374 562226
rect 435430 562170 435498 562226
rect 435554 562170 435622 562226
rect 435678 562170 435774 562226
rect 435154 562102 435774 562170
rect 435154 562046 435250 562102
rect 435306 562046 435374 562102
rect 435430 562046 435498 562102
rect 435554 562046 435622 562102
rect 435678 562046 435774 562102
rect 435154 561978 435774 562046
rect 435154 561922 435250 561978
rect 435306 561922 435374 561978
rect 435430 561922 435498 561978
rect 435554 561922 435622 561978
rect 435678 561922 435774 561978
rect 435154 544350 435774 561922
rect 435154 544294 435250 544350
rect 435306 544294 435374 544350
rect 435430 544294 435498 544350
rect 435554 544294 435622 544350
rect 435678 544294 435774 544350
rect 435154 544226 435774 544294
rect 435154 544170 435250 544226
rect 435306 544170 435374 544226
rect 435430 544170 435498 544226
rect 435554 544170 435622 544226
rect 435678 544170 435774 544226
rect 435154 544102 435774 544170
rect 435154 544046 435250 544102
rect 435306 544046 435374 544102
rect 435430 544046 435498 544102
rect 435554 544046 435622 544102
rect 435678 544046 435774 544102
rect 435154 543978 435774 544046
rect 435154 543922 435250 543978
rect 435306 543922 435374 543978
rect 435430 543922 435498 543978
rect 435554 543922 435622 543978
rect 435678 543922 435774 543978
rect 435154 527750 435774 543922
rect 438874 598172 439494 598268
rect 438874 598116 438970 598172
rect 439026 598116 439094 598172
rect 439150 598116 439218 598172
rect 439274 598116 439342 598172
rect 439398 598116 439494 598172
rect 438874 598048 439494 598116
rect 438874 597992 438970 598048
rect 439026 597992 439094 598048
rect 439150 597992 439218 598048
rect 439274 597992 439342 598048
rect 439398 597992 439494 598048
rect 438874 597924 439494 597992
rect 438874 597868 438970 597924
rect 439026 597868 439094 597924
rect 439150 597868 439218 597924
rect 439274 597868 439342 597924
rect 439398 597868 439494 597924
rect 438874 597800 439494 597868
rect 438874 597744 438970 597800
rect 439026 597744 439094 597800
rect 439150 597744 439218 597800
rect 439274 597744 439342 597800
rect 439398 597744 439494 597800
rect 438874 586350 439494 597744
rect 438874 586294 438970 586350
rect 439026 586294 439094 586350
rect 439150 586294 439218 586350
rect 439274 586294 439342 586350
rect 439398 586294 439494 586350
rect 438874 586226 439494 586294
rect 438874 586170 438970 586226
rect 439026 586170 439094 586226
rect 439150 586170 439218 586226
rect 439274 586170 439342 586226
rect 439398 586170 439494 586226
rect 438874 586102 439494 586170
rect 438874 586046 438970 586102
rect 439026 586046 439094 586102
rect 439150 586046 439218 586102
rect 439274 586046 439342 586102
rect 439398 586046 439494 586102
rect 438874 585978 439494 586046
rect 438874 585922 438970 585978
rect 439026 585922 439094 585978
rect 439150 585922 439218 585978
rect 439274 585922 439342 585978
rect 439398 585922 439494 585978
rect 438874 568350 439494 585922
rect 438874 568294 438970 568350
rect 439026 568294 439094 568350
rect 439150 568294 439218 568350
rect 439274 568294 439342 568350
rect 439398 568294 439494 568350
rect 438874 568226 439494 568294
rect 438874 568170 438970 568226
rect 439026 568170 439094 568226
rect 439150 568170 439218 568226
rect 439274 568170 439342 568226
rect 439398 568170 439494 568226
rect 438874 568102 439494 568170
rect 438874 568046 438970 568102
rect 439026 568046 439094 568102
rect 439150 568046 439218 568102
rect 439274 568046 439342 568102
rect 439398 568046 439494 568102
rect 438874 567978 439494 568046
rect 438874 567922 438970 567978
rect 439026 567922 439094 567978
rect 439150 567922 439218 567978
rect 439274 567922 439342 567978
rect 439398 567922 439494 567978
rect 438874 550350 439494 567922
rect 438874 550294 438970 550350
rect 439026 550294 439094 550350
rect 439150 550294 439218 550350
rect 439274 550294 439342 550350
rect 439398 550294 439494 550350
rect 438874 550226 439494 550294
rect 438874 550170 438970 550226
rect 439026 550170 439094 550226
rect 439150 550170 439218 550226
rect 439274 550170 439342 550226
rect 439398 550170 439494 550226
rect 438874 550102 439494 550170
rect 438874 550046 438970 550102
rect 439026 550046 439094 550102
rect 439150 550046 439218 550102
rect 439274 550046 439342 550102
rect 439398 550046 439494 550102
rect 438874 549978 439494 550046
rect 438874 549922 438970 549978
rect 439026 549922 439094 549978
rect 439150 549922 439218 549978
rect 439274 549922 439342 549978
rect 439398 549922 439494 549978
rect 438874 532350 439494 549922
rect 438874 532294 438970 532350
rect 439026 532294 439094 532350
rect 439150 532294 439218 532350
rect 439274 532294 439342 532350
rect 439398 532294 439494 532350
rect 438874 532226 439494 532294
rect 438874 532170 438970 532226
rect 439026 532170 439094 532226
rect 439150 532170 439218 532226
rect 439274 532170 439342 532226
rect 439398 532170 439494 532226
rect 438874 532102 439494 532170
rect 438874 532046 438970 532102
rect 439026 532046 439094 532102
rect 439150 532046 439218 532102
rect 439274 532046 439342 532102
rect 439398 532046 439494 532102
rect 438874 531978 439494 532046
rect 438874 531922 438970 531978
rect 439026 531922 439094 531978
rect 439150 531922 439218 531978
rect 439274 531922 439342 531978
rect 439398 531922 439494 531978
rect 438874 527750 439494 531922
rect 453154 597212 453774 598268
rect 453154 597156 453250 597212
rect 453306 597156 453374 597212
rect 453430 597156 453498 597212
rect 453554 597156 453622 597212
rect 453678 597156 453774 597212
rect 453154 597088 453774 597156
rect 453154 597032 453250 597088
rect 453306 597032 453374 597088
rect 453430 597032 453498 597088
rect 453554 597032 453622 597088
rect 453678 597032 453774 597088
rect 453154 596964 453774 597032
rect 453154 596908 453250 596964
rect 453306 596908 453374 596964
rect 453430 596908 453498 596964
rect 453554 596908 453622 596964
rect 453678 596908 453774 596964
rect 453154 596840 453774 596908
rect 453154 596784 453250 596840
rect 453306 596784 453374 596840
rect 453430 596784 453498 596840
rect 453554 596784 453622 596840
rect 453678 596784 453774 596840
rect 453154 580350 453774 596784
rect 453154 580294 453250 580350
rect 453306 580294 453374 580350
rect 453430 580294 453498 580350
rect 453554 580294 453622 580350
rect 453678 580294 453774 580350
rect 453154 580226 453774 580294
rect 453154 580170 453250 580226
rect 453306 580170 453374 580226
rect 453430 580170 453498 580226
rect 453554 580170 453622 580226
rect 453678 580170 453774 580226
rect 453154 580102 453774 580170
rect 453154 580046 453250 580102
rect 453306 580046 453374 580102
rect 453430 580046 453498 580102
rect 453554 580046 453622 580102
rect 453678 580046 453774 580102
rect 453154 579978 453774 580046
rect 453154 579922 453250 579978
rect 453306 579922 453374 579978
rect 453430 579922 453498 579978
rect 453554 579922 453622 579978
rect 453678 579922 453774 579978
rect 453154 562350 453774 579922
rect 453154 562294 453250 562350
rect 453306 562294 453374 562350
rect 453430 562294 453498 562350
rect 453554 562294 453622 562350
rect 453678 562294 453774 562350
rect 453154 562226 453774 562294
rect 453154 562170 453250 562226
rect 453306 562170 453374 562226
rect 453430 562170 453498 562226
rect 453554 562170 453622 562226
rect 453678 562170 453774 562226
rect 453154 562102 453774 562170
rect 453154 562046 453250 562102
rect 453306 562046 453374 562102
rect 453430 562046 453498 562102
rect 453554 562046 453622 562102
rect 453678 562046 453774 562102
rect 453154 561978 453774 562046
rect 453154 561922 453250 561978
rect 453306 561922 453374 561978
rect 453430 561922 453498 561978
rect 453554 561922 453622 561978
rect 453678 561922 453774 561978
rect 453154 544350 453774 561922
rect 453154 544294 453250 544350
rect 453306 544294 453374 544350
rect 453430 544294 453498 544350
rect 453554 544294 453622 544350
rect 453678 544294 453774 544350
rect 453154 544226 453774 544294
rect 453154 544170 453250 544226
rect 453306 544170 453374 544226
rect 453430 544170 453498 544226
rect 453554 544170 453622 544226
rect 453678 544170 453774 544226
rect 453154 544102 453774 544170
rect 453154 544046 453250 544102
rect 453306 544046 453374 544102
rect 453430 544046 453498 544102
rect 453554 544046 453622 544102
rect 453678 544046 453774 544102
rect 453154 543978 453774 544046
rect 453154 543922 453250 543978
rect 453306 543922 453374 543978
rect 453430 543922 453498 543978
rect 453554 543922 453622 543978
rect 453678 543922 453774 543978
rect 453154 528388 453774 543922
rect 456874 598172 457494 598268
rect 456874 598116 456970 598172
rect 457026 598116 457094 598172
rect 457150 598116 457218 598172
rect 457274 598116 457342 598172
rect 457398 598116 457494 598172
rect 456874 598048 457494 598116
rect 456874 597992 456970 598048
rect 457026 597992 457094 598048
rect 457150 597992 457218 598048
rect 457274 597992 457342 598048
rect 457398 597992 457494 598048
rect 456874 597924 457494 597992
rect 456874 597868 456970 597924
rect 457026 597868 457094 597924
rect 457150 597868 457218 597924
rect 457274 597868 457342 597924
rect 457398 597868 457494 597924
rect 456874 597800 457494 597868
rect 456874 597744 456970 597800
rect 457026 597744 457094 597800
rect 457150 597744 457218 597800
rect 457274 597744 457342 597800
rect 457398 597744 457494 597800
rect 456874 586350 457494 597744
rect 456874 586294 456970 586350
rect 457026 586294 457094 586350
rect 457150 586294 457218 586350
rect 457274 586294 457342 586350
rect 457398 586294 457494 586350
rect 456874 586226 457494 586294
rect 456874 586170 456970 586226
rect 457026 586170 457094 586226
rect 457150 586170 457218 586226
rect 457274 586170 457342 586226
rect 457398 586170 457494 586226
rect 456874 586102 457494 586170
rect 456874 586046 456970 586102
rect 457026 586046 457094 586102
rect 457150 586046 457218 586102
rect 457274 586046 457342 586102
rect 457398 586046 457494 586102
rect 456874 585978 457494 586046
rect 456874 585922 456970 585978
rect 457026 585922 457094 585978
rect 457150 585922 457218 585978
rect 457274 585922 457342 585978
rect 457398 585922 457494 585978
rect 456874 568350 457494 585922
rect 456874 568294 456970 568350
rect 457026 568294 457094 568350
rect 457150 568294 457218 568350
rect 457274 568294 457342 568350
rect 457398 568294 457494 568350
rect 456874 568226 457494 568294
rect 456874 568170 456970 568226
rect 457026 568170 457094 568226
rect 457150 568170 457218 568226
rect 457274 568170 457342 568226
rect 457398 568170 457494 568226
rect 456874 568102 457494 568170
rect 456874 568046 456970 568102
rect 457026 568046 457094 568102
rect 457150 568046 457218 568102
rect 457274 568046 457342 568102
rect 457398 568046 457494 568102
rect 456874 567978 457494 568046
rect 456874 567922 456970 567978
rect 457026 567922 457094 567978
rect 457150 567922 457218 567978
rect 457274 567922 457342 567978
rect 457398 567922 457494 567978
rect 456874 550350 457494 567922
rect 456874 550294 456970 550350
rect 457026 550294 457094 550350
rect 457150 550294 457218 550350
rect 457274 550294 457342 550350
rect 457398 550294 457494 550350
rect 456874 550226 457494 550294
rect 456874 550170 456970 550226
rect 457026 550170 457094 550226
rect 457150 550170 457218 550226
rect 457274 550170 457342 550226
rect 457398 550170 457494 550226
rect 456874 550102 457494 550170
rect 456874 550046 456970 550102
rect 457026 550046 457094 550102
rect 457150 550046 457218 550102
rect 457274 550046 457342 550102
rect 457398 550046 457494 550102
rect 456874 549978 457494 550046
rect 456874 549922 456970 549978
rect 457026 549922 457094 549978
rect 457150 549922 457218 549978
rect 457274 549922 457342 549978
rect 457398 549922 457494 549978
rect 456874 532350 457494 549922
rect 456874 532294 456970 532350
rect 457026 532294 457094 532350
rect 457150 532294 457218 532350
rect 457274 532294 457342 532350
rect 457398 532294 457494 532350
rect 456874 532226 457494 532294
rect 456874 532170 456970 532226
rect 457026 532170 457094 532226
rect 457150 532170 457218 532226
rect 457274 532170 457342 532226
rect 457398 532170 457494 532226
rect 456874 532102 457494 532170
rect 456874 532046 456970 532102
rect 457026 532046 457094 532102
rect 457150 532046 457218 532102
rect 457274 532046 457342 532102
rect 457398 532046 457494 532102
rect 456874 531978 457494 532046
rect 456874 531922 456970 531978
rect 457026 531922 457094 531978
rect 457150 531922 457218 531978
rect 457274 531922 457342 531978
rect 457398 531922 457494 531978
rect 456874 527750 457494 531922
rect 471154 597212 471774 598268
rect 471154 597156 471250 597212
rect 471306 597156 471374 597212
rect 471430 597156 471498 597212
rect 471554 597156 471622 597212
rect 471678 597156 471774 597212
rect 471154 597088 471774 597156
rect 471154 597032 471250 597088
rect 471306 597032 471374 597088
rect 471430 597032 471498 597088
rect 471554 597032 471622 597088
rect 471678 597032 471774 597088
rect 471154 596964 471774 597032
rect 471154 596908 471250 596964
rect 471306 596908 471374 596964
rect 471430 596908 471498 596964
rect 471554 596908 471622 596964
rect 471678 596908 471774 596964
rect 471154 596840 471774 596908
rect 471154 596784 471250 596840
rect 471306 596784 471374 596840
rect 471430 596784 471498 596840
rect 471554 596784 471622 596840
rect 471678 596784 471774 596840
rect 471154 580350 471774 596784
rect 471154 580294 471250 580350
rect 471306 580294 471374 580350
rect 471430 580294 471498 580350
rect 471554 580294 471622 580350
rect 471678 580294 471774 580350
rect 471154 580226 471774 580294
rect 471154 580170 471250 580226
rect 471306 580170 471374 580226
rect 471430 580170 471498 580226
rect 471554 580170 471622 580226
rect 471678 580170 471774 580226
rect 471154 580102 471774 580170
rect 471154 580046 471250 580102
rect 471306 580046 471374 580102
rect 471430 580046 471498 580102
rect 471554 580046 471622 580102
rect 471678 580046 471774 580102
rect 471154 579978 471774 580046
rect 471154 579922 471250 579978
rect 471306 579922 471374 579978
rect 471430 579922 471498 579978
rect 471554 579922 471622 579978
rect 471678 579922 471774 579978
rect 471154 562350 471774 579922
rect 471154 562294 471250 562350
rect 471306 562294 471374 562350
rect 471430 562294 471498 562350
rect 471554 562294 471622 562350
rect 471678 562294 471774 562350
rect 471154 562226 471774 562294
rect 471154 562170 471250 562226
rect 471306 562170 471374 562226
rect 471430 562170 471498 562226
rect 471554 562170 471622 562226
rect 471678 562170 471774 562226
rect 471154 562102 471774 562170
rect 471154 562046 471250 562102
rect 471306 562046 471374 562102
rect 471430 562046 471498 562102
rect 471554 562046 471622 562102
rect 471678 562046 471774 562102
rect 471154 561978 471774 562046
rect 471154 561922 471250 561978
rect 471306 561922 471374 561978
rect 471430 561922 471498 561978
rect 471554 561922 471622 561978
rect 471678 561922 471774 561978
rect 471154 544350 471774 561922
rect 471154 544294 471250 544350
rect 471306 544294 471374 544350
rect 471430 544294 471498 544350
rect 471554 544294 471622 544350
rect 471678 544294 471774 544350
rect 471154 544226 471774 544294
rect 471154 544170 471250 544226
rect 471306 544170 471374 544226
rect 471430 544170 471498 544226
rect 471554 544170 471622 544226
rect 471678 544170 471774 544226
rect 471154 544102 471774 544170
rect 471154 544046 471250 544102
rect 471306 544046 471374 544102
rect 471430 544046 471498 544102
rect 471554 544046 471622 544102
rect 471678 544046 471774 544102
rect 471154 543978 471774 544046
rect 471154 543922 471250 543978
rect 471306 543922 471374 543978
rect 471430 543922 471498 543978
rect 471554 543922 471622 543978
rect 471678 543922 471774 543978
rect 471154 527750 471774 543922
rect 474874 598172 475494 598268
rect 474874 598116 474970 598172
rect 475026 598116 475094 598172
rect 475150 598116 475218 598172
rect 475274 598116 475342 598172
rect 475398 598116 475494 598172
rect 474874 598048 475494 598116
rect 474874 597992 474970 598048
rect 475026 597992 475094 598048
rect 475150 597992 475218 598048
rect 475274 597992 475342 598048
rect 475398 597992 475494 598048
rect 474874 597924 475494 597992
rect 474874 597868 474970 597924
rect 475026 597868 475094 597924
rect 475150 597868 475218 597924
rect 475274 597868 475342 597924
rect 475398 597868 475494 597924
rect 474874 597800 475494 597868
rect 474874 597744 474970 597800
rect 475026 597744 475094 597800
rect 475150 597744 475218 597800
rect 475274 597744 475342 597800
rect 475398 597744 475494 597800
rect 474874 586350 475494 597744
rect 474874 586294 474970 586350
rect 475026 586294 475094 586350
rect 475150 586294 475218 586350
rect 475274 586294 475342 586350
rect 475398 586294 475494 586350
rect 474874 586226 475494 586294
rect 474874 586170 474970 586226
rect 475026 586170 475094 586226
rect 475150 586170 475218 586226
rect 475274 586170 475342 586226
rect 475398 586170 475494 586226
rect 474874 586102 475494 586170
rect 474874 586046 474970 586102
rect 475026 586046 475094 586102
rect 475150 586046 475218 586102
rect 475274 586046 475342 586102
rect 475398 586046 475494 586102
rect 474874 585978 475494 586046
rect 474874 585922 474970 585978
rect 475026 585922 475094 585978
rect 475150 585922 475218 585978
rect 475274 585922 475342 585978
rect 475398 585922 475494 585978
rect 474874 568350 475494 585922
rect 474874 568294 474970 568350
rect 475026 568294 475094 568350
rect 475150 568294 475218 568350
rect 475274 568294 475342 568350
rect 475398 568294 475494 568350
rect 474874 568226 475494 568294
rect 474874 568170 474970 568226
rect 475026 568170 475094 568226
rect 475150 568170 475218 568226
rect 475274 568170 475342 568226
rect 475398 568170 475494 568226
rect 474874 568102 475494 568170
rect 474874 568046 474970 568102
rect 475026 568046 475094 568102
rect 475150 568046 475218 568102
rect 475274 568046 475342 568102
rect 475398 568046 475494 568102
rect 474874 567978 475494 568046
rect 474874 567922 474970 567978
rect 475026 567922 475094 567978
rect 475150 567922 475218 567978
rect 475274 567922 475342 567978
rect 475398 567922 475494 567978
rect 474874 550350 475494 567922
rect 474874 550294 474970 550350
rect 475026 550294 475094 550350
rect 475150 550294 475218 550350
rect 475274 550294 475342 550350
rect 475398 550294 475494 550350
rect 474874 550226 475494 550294
rect 474874 550170 474970 550226
rect 475026 550170 475094 550226
rect 475150 550170 475218 550226
rect 475274 550170 475342 550226
rect 475398 550170 475494 550226
rect 474874 550102 475494 550170
rect 474874 550046 474970 550102
rect 475026 550046 475094 550102
rect 475150 550046 475218 550102
rect 475274 550046 475342 550102
rect 475398 550046 475494 550102
rect 474874 549978 475494 550046
rect 474874 549922 474970 549978
rect 475026 549922 475094 549978
rect 475150 549922 475218 549978
rect 475274 549922 475342 549978
rect 475398 549922 475494 549978
rect 474874 532350 475494 549922
rect 474874 532294 474970 532350
rect 475026 532294 475094 532350
rect 475150 532294 475218 532350
rect 475274 532294 475342 532350
rect 475398 532294 475494 532350
rect 474874 532226 475494 532294
rect 474874 532170 474970 532226
rect 475026 532170 475094 532226
rect 475150 532170 475218 532226
rect 475274 532170 475342 532226
rect 475398 532170 475494 532226
rect 474874 532102 475494 532170
rect 474874 532046 474970 532102
rect 475026 532046 475094 532102
rect 475150 532046 475218 532102
rect 475274 532046 475342 532102
rect 475398 532046 475494 532102
rect 474874 531978 475494 532046
rect 474874 531922 474970 531978
rect 475026 531922 475094 531978
rect 475150 531922 475218 531978
rect 475274 531922 475342 531978
rect 475398 531922 475494 531978
rect 474874 527750 475494 531922
rect 489154 597212 489774 598268
rect 489154 597156 489250 597212
rect 489306 597156 489374 597212
rect 489430 597156 489498 597212
rect 489554 597156 489622 597212
rect 489678 597156 489774 597212
rect 489154 597088 489774 597156
rect 489154 597032 489250 597088
rect 489306 597032 489374 597088
rect 489430 597032 489498 597088
rect 489554 597032 489622 597088
rect 489678 597032 489774 597088
rect 489154 596964 489774 597032
rect 489154 596908 489250 596964
rect 489306 596908 489374 596964
rect 489430 596908 489498 596964
rect 489554 596908 489622 596964
rect 489678 596908 489774 596964
rect 489154 596840 489774 596908
rect 489154 596784 489250 596840
rect 489306 596784 489374 596840
rect 489430 596784 489498 596840
rect 489554 596784 489622 596840
rect 489678 596784 489774 596840
rect 489154 580350 489774 596784
rect 489154 580294 489250 580350
rect 489306 580294 489374 580350
rect 489430 580294 489498 580350
rect 489554 580294 489622 580350
rect 489678 580294 489774 580350
rect 489154 580226 489774 580294
rect 489154 580170 489250 580226
rect 489306 580170 489374 580226
rect 489430 580170 489498 580226
rect 489554 580170 489622 580226
rect 489678 580170 489774 580226
rect 489154 580102 489774 580170
rect 489154 580046 489250 580102
rect 489306 580046 489374 580102
rect 489430 580046 489498 580102
rect 489554 580046 489622 580102
rect 489678 580046 489774 580102
rect 489154 579978 489774 580046
rect 489154 579922 489250 579978
rect 489306 579922 489374 579978
rect 489430 579922 489498 579978
rect 489554 579922 489622 579978
rect 489678 579922 489774 579978
rect 489154 562350 489774 579922
rect 489154 562294 489250 562350
rect 489306 562294 489374 562350
rect 489430 562294 489498 562350
rect 489554 562294 489622 562350
rect 489678 562294 489774 562350
rect 489154 562226 489774 562294
rect 489154 562170 489250 562226
rect 489306 562170 489374 562226
rect 489430 562170 489498 562226
rect 489554 562170 489622 562226
rect 489678 562170 489774 562226
rect 489154 562102 489774 562170
rect 489154 562046 489250 562102
rect 489306 562046 489374 562102
rect 489430 562046 489498 562102
rect 489554 562046 489622 562102
rect 489678 562046 489774 562102
rect 489154 561978 489774 562046
rect 489154 561922 489250 561978
rect 489306 561922 489374 561978
rect 489430 561922 489498 561978
rect 489554 561922 489622 561978
rect 489678 561922 489774 561978
rect 489154 544350 489774 561922
rect 489154 544294 489250 544350
rect 489306 544294 489374 544350
rect 489430 544294 489498 544350
rect 489554 544294 489622 544350
rect 489678 544294 489774 544350
rect 489154 544226 489774 544294
rect 489154 544170 489250 544226
rect 489306 544170 489374 544226
rect 489430 544170 489498 544226
rect 489554 544170 489622 544226
rect 489678 544170 489774 544226
rect 489154 544102 489774 544170
rect 489154 544046 489250 544102
rect 489306 544046 489374 544102
rect 489430 544046 489498 544102
rect 489554 544046 489622 544102
rect 489678 544046 489774 544102
rect 489154 543978 489774 544046
rect 489154 543922 489250 543978
rect 489306 543922 489374 543978
rect 489430 543922 489498 543978
rect 489554 543922 489622 543978
rect 489678 543922 489774 543978
rect 489154 527750 489774 543922
rect 492874 598172 493494 598268
rect 492874 598116 492970 598172
rect 493026 598116 493094 598172
rect 493150 598116 493218 598172
rect 493274 598116 493342 598172
rect 493398 598116 493494 598172
rect 492874 598048 493494 598116
rect 492874 597992 492970 598048
rect 493026 597992 493094 598048
rect 493150 597992 493218 598048
rect 493274 597992 493342 598048
rect 493398 597992 493494 598048
rect 492874 597924 493494 597992
rect 492874 597868 492970 597924
rect 493026 597868 493094 597924
rect 493150 597868 493218 597924
rect 493274 597868 493342 597924
rect 493398 597868 493494 597924
rect 492874 597800 493494 597868
rect 492874 597744 492970 597800
rect 493026 597744 493094 597800
rect 493150 597744 493218 597800
rect 493274 597744 493342 597800
rect 493398 597744 493494 597800
rect 492874 586350 493494 597744
rect 492874 586294 492970 586350
rect 493026 586294 493094 586350
rect 493150 586294 493218 586350
rect 493274 586294 493342 586350
rect 493398 586294 493494 586350
rect 492874 586226 493494 586294
rect 492874 586170 492970 586226
rect 493026 586170 493094 586226
rect 493150 586170 493218 586226
rect 493274 586170 493342 586226
rect 493398 586170 493494 586226
rect 492874 586102 493494 586170
rect 492874 586046 492970 586102
rect 493026 586046 493094 586102
rect 493150 586046 493218 586102
rect 493274 586046 493342 586102
rect 493398 586046 493494 586102
rect 492874 585978 493494 586046
rect 492874 585922 492970 585978
rect 493026 585922 493094 585978
rect 493150 585922 493218 585978
rect 493274 585922 493342 585978
rect 493398 585922 493494 585978
rect 492874 568350 493494 585922
rect 492874 568294 492970 568350
rect 493026 568294 493094 568350
rect 493150 568294 493218 568350
rect 493274 568294 493342 568350
rect 493398 568294 493494 568350
rect 492874 568226 493494 568294
rect 492874 568170 492970 568226
rect 493026 568170 493094 568226
rect 493150 568170 493218 568226
rect 493274 568170 493342 568226
rect 493398 568170 493494 568226
rect 492874 568102 493494 568170
rect 492874 568046 492970 568102
rect 493026 568046 493094 568102
rect 493150 568046 493218 568102
rect 493274 568046 493342 568102
rect 493398 568046 493494 568102
rect 492874 567978 493494 568046
rect 492874 567922 492970 567978
rect 493026 567922 493094 567978
rect 493150 567922 493218 567978
rect 493274 567922 493342 567978
rect 493398 567922 493494 567978
rect 492874 550350 493494 567922
rect 492874 550294 492970 550350
rect 493026 550294 493094 550350
rect 493150 550294 493218 550350
rect 493274 550294 493342 550350
rect 493398 550294 493494 550350
rect 492874 550226 493494 550294
rect 492874 550170 492970 550226
rect 493026 550170 493094 550226
rect 493150 550170 493218 550226
rect 493274 550170 493342 550226
rect 493398 550170 493494 550226
rect 492874 550102 493494 550170
rect 492874 550046 492970 550102
rect 493026 550046 493094 550102
rect 493150 550046 493218 550102
rect 493274 550046 493342 550102
rect 493398 550046 493494 550102
rect 492874 549978 493494 550046
rect 492874 549922 492970 549978
rect 493026 549922 493094 549978
rect 493150 549922 493218 549978
rect 493274 549922 493342 549978
rect 493398 549922 493494 549978
rect 492874 532350 493494 549922
rect 492874 532294 492970 532350
rect 493026 532294 493094 532350
rect 493150 532294 493218 532350
rect 493274 532294 493342 532350
rect 493398 532294 493494 532350
rect 492874 532226 493494 532294
rect 492874 532170 492970 532226
rect 493026 532170 493094 532226
rect 493150 532170 493218 532226
rect 493274 532170 493342 532226
rect 493398 532170 493494 532226
rect 492874 532102 493494 532170
rect 492874 532046 492970 532102
rect 493026 532046 493094 532102
rect 493150 532046 493218 532102
rect 493274 532046 493342 532102
rect 493398 532046 493494 532102
rect 492874 531978 493494 532046
rect 492874 531922 492970 531978
rect 493026 531922 493094 531978
rect 493150 531922 493218 531978
rect 493274 531922 493342 531978
rect 493398 531922 493494 531978
rect 492874 527750 493494 531922
rect 507154 597212 507774 598268
rect 507154 597156 507250 597212
rect 507306 597156 507374 597212
rect 507430 597156 507498 597212
rect 507554 597156 507622 597212
rect 507678 597156 507774 597212
rect 507154 597088 507774 597156
rect 507154 597032 507250 597088
rect 507306 597032 507374 597088
rect 507430 597032 507498 597088
rect 507554 597032 507622 597088
rect 507678 597032 507774 597088
rect 507154 596964 507774 597032
rect 507154 596908 507250 596964
rect 507306 596908 507374 596964
rect 507430 596908 507498 596964
rect 507554 596908 507622 596964
rect 507678 596908 507774 596964
rect 507154 596840 507774 596908
rect 507154 596784 507250 596840
rect 507306 596784 507374 596840
rect 507430 596784 507498 596840
rect 507554 596784 507622 596840
rect 507678 596784 507774 596840
rect 507154 580350 507774 596784
rect 507154 580294 507250 580350
rect 507306 580294 507374 580350
rect 507430 580294 507498 580350
rect 507554 580294 507622 580350
rect 507678 580294 507774 580350
rect 507154 580226 507774 580294
rect 507154 580170 507250 580226
rect 507306 580170 507374 580226
rect 507430 580170 507498 580226
rect 507554 580170 507622 580226
rect 507678 580170 507774 580226
rect 507154 580102 507774 580170
rect 507154 580046 507250 580102
rect 507306 580046 507374 580102
rect 507430 580046 507498 580102
rect 507554 580046 507622 580102
rect 507678 580046 507774 580102
rect 507154 579978 507774 580046
rect 507154 579922 507250 579978
rect 507306 579922 507374 579978
rect 507430 579922 507498 579978
rect 507554 579922 507622 579978
rect 507678 579922 507774 579978
rect 507154 562350 507774 579922
rect 507154 562294 507250 562350
rect 507306 562294 507374 562350
rect 507430 562294 507498 562350
rect 507554 562294 507622 562350
rect 507678 562294 507774 562350
rect 507154 562226 507774 562294
rect 507154 562170 507250 562226
rect 507306 562170 507374 562226
rect 507430 562170 507498 562226
rect 507554 562170 507622 562226
rect 507678 562170 507774 562226
rect 507154 562102 507774 562170
rect 507154 562046 507250 562102
rect 507306 562046 507374 562102
rect 507430 562046 507498 562102
rect 507554 562046 507622 562102
rect 507678 562046 507774 562102
rect 507154 561978 507774 562046
rect 507154 561922 507250 561978
rect 507306 561922 507374 561978
rect 507430 561922 507498 561978
rect 507554 561922 507622 561978
rect 507678 561922 507774 561978
rect 507154 544350 507774 561922
rect 507154 544294 507250 544350
rect 507306 544294 507374 544350
rect 507430 544294 507498 544350
rect 507554 544294 507622 544350
rect 507678 544294 507774 544350
rect 507154 544226 507774 544294
rect 507154 544170 507250 544226
rect 507306 544170 507374 544226
rect 507430 544170 507498 544226
rect 507554 544170 507622 544226
rect 507678 544170 507774 544226
rect 507154 544102 507774 544170
rect 507154 544046 507250 544102
rect 507306 544046 507374 544102
rect 507430 544046 507498 544102
rect 507554 544046 507622 544102
rect 507678 544046 507774 544102
rect 507154 543978 507774 544046
rect 507154 543922 507250 543978
rect 507306 543922 507374 543978
rect 507430 543922 507498 543978
rect 507554 543922 507622 543978
rect 507678 543922 507774 543978
rect 507154 527750 507774 543922
rect 510874 598172 511494 598268
rect 510874 598116 510970 598172
rect 511026 598116 511094 598172
rect 511150 598116 511218 598172
rect 511274 598116 511342 598172
rect 511398 598116 511494 598172
rect 510874 598048 511494 598116
rect 510874 597992 510970 598048
rect 511026 597992 511094 598048
rect 511150 597992 511218 598048
rect 511274 597992 511342 598048
rect 511398 597992 511494 598048
rect 510874 597924 511494 597992
rect 510874 597868 510970 597924
rect 511026 597868 511094 597924
rect 511150 597868 511218 597924
rect 511274 597868 511342 597924
rect 511398 597868 511494 597924
rect 510874 597800 511494 597868
rect 510874 597744 510970 597800
rect 511026 597744 511094 597800
rect 511150 597744 511218 597800
rect 511274 597744 511342 597800
rect 511398 597744 511494 597800
rect 510874 586350 511494 597744
rect 510874 586294 510970 586350
rect 511026 586294 511094 586350
rect 511150 586294 511218 586350
rect 511274 586294 511342 586350
rect 511398 586294 511494 586350
rect 510874 586226 511494 586294
rect 510874 586170 510970 586226
rect 511026 586170 511094 586226
rect 511150 586170 511218 586226
rect 511274 586170 511342 586226
rect 511398 586170 511494 586226
rect 510874 586102 511494 586170
rect 510874 586046 510970 586102
rect 511026 586046 511094 586102
rect 511150 586046 511218 586102
rect 511274 586046 511342 586102
rect 511398 586046 511494 586102
rect 510874 585978 511494 586046
rect 510874 585922 510970 585978
rect 511026 585922 511094 585978
rect 511150 585922 511218 585978
rect 511274 585922 511342 585978
rect 511398 585922 511494 585978
rect 510874 568350 511494 585922
rect 510874 568294 510970 568350
rect 511026 568294 511094 568350
rect 511150 568294 511218 568350
rect 511274 568294 511342 568350
rect 511398 568294 511494 568350
rect 510874 568226 511494 568294
rect 510874 568170 510970 568226
rect 511026 568170 511094 568226
rect 511150 568170 511218 568226
rect 511274 568170 511342 568226
rect 511398 568170 511494 568226
rect 510874 568102 511494 568170
rect 510874 568046 510970 568102
rect 511026 568046 511094 568102
rect 511150 568046 511218 568102
rect 511274 568046 511342 568102
rect 511398 568046 511494 568102
rect 510874 567978 511494 568046
rect 510874 567922 510970 567978
rect 511026 567922 511094 567978
rect 511150 567922 511218 567978
rect 511274 567922 511342 567978
rect 511398 567922 511494 567978
rect 510874 550350 511494 567922
rect 510874 550294 510970 550350
rect 511026 550294 511094 550350
rect 511150 550294 511218 550350
rect 511274 550294 511342 550350
rect 511398 550294 511494 550350
rect 510874 550226 511494 550294
rect 510874 550170 510970 550226
rect 511026 550170 511094 550226
rect 511150 550170 511218 550226
rect 511274 550170 511342 550226
rect 511398 550170 511494 550226
rect 510874 550102 511494 550170
rect 510874 550046 510970 550102
rect 511026 550046 511094 550102
rect 511150 550046 511218 550102
rect 511274 550046 511342 550102
rect 511398 550046 511494 550102
rect 510874 549978 511494 550046
rect 510874 549922 510970 549978
rect 511026 549922 511094 549978
rect 511150 549922 511218 549978
rect 511274 549922 511342 549978
rect 511398 549922 511494 549978
rect 510874 532350 511494 549922
rect 510874 532294 510970 532350
rect 511026 532294 511094 532350
rect 511150 532294 511218 532350
rect 511274 532294 511342 532350
rect 511398 532294 511494 532350
rect 510874 532226 511494 532294
rect 510874 532170 510970 532226
rect 511026 532170 511094 532226
rect 511150 532170 511218 532226
rect 511274 532170 511342 532226
rect 511398 532170 511494 532226
rect 510874 532102 511494 532170
rect 510874 532046 510970 532102
rect 511026 532046 511094 532102
rect 511150 532046 511218 532102
rect 511274 532046 511342 532102
rect 511398 532046 511494 532102
rect 510874 531978 511494 532046
rect 510874 531922 510970 531978
rect 511026 531922 511094 531978
rect 511150 531922 511218 531978
rect 511274 531922 511342 531978
rect 511398 531922 511494 531978
rect 510874 527750 511494 531922
rect 525154 597212 525774 598268
rect 525154 597156 525250 597212
rect 525306 597156 525374 597212
rect 525430 597156 525498 597212
rect 525554 597156 525622 597212
rect 525678 597156 525774 597212
rect 525154 597088 525774 597156
rect 525154 597032 525250 597088
rect 525306 597032 525374 597088
rect 525430 597032 525498 597088
rect 525554 597032 525622 597088
rect 525678 597032 525774 597088
rect 525154 596964 525774 597032
rect 525154 596908 525250 596964
rect 525306 596908 525374 596964
rect 525430 596908 525498 596964
rect 525554 596908 525622 596964
rect 525678 596908 525774 596964
rect 525154 596840 525774 596908
rect 525154 596784 525250 596840
rect 525306 596784 525374 596840
rect 525430 596784 525498 596840
rect 525554 596784 525622 596840
rect 525678 596784 525774 596840
rect 525154 580350 525774 596784
rect 525154 580294 525250 580350
rect 525306 580294 525374 580350
rect 525430 580294 525498 580350
rect 525554 580294 525622 580350
rect 525678 580294 525774 580350
rect 525154 580226 525774 580294
rect 525154 580170 525250 580226
rect 525306 580170 525374 580226
rect 525430 580170 525498 580226
rect 525554 580170 525622 580226
rect 525678 580170 525774 580226
rect 525154 580102 525774 580170
rect 525154 580046 525250 580102
rect 525306 580046 525374 580102
rect 525430 580046 525498 580102
rect 525554 580046 525622 580102
rect 525678 580046 525774 580102
rect 525154 579978 525774 580046
rect 525154 579922 525250 579978
rect 525306 579922 525374 579978
rect 525430 579922 525498 579978
rect 525554 579922 525622 579978
rect 525678 579922 525774 579978
rect 525154 562350 525774 579922
rect 525154 562294 525250 562350
rect 525306 562294 525374 562350
rect 525430 562294 525498 562350
rect 525554 562294 525622 562350
rect 525678 562294 525774 562350
rect 525154 562226 525774 562294
rect 525154 562170 525250 562226
rect 525306 562170 525374 562226
rect 525430 562170 525498 562226
rect 525554 562170 525622 562226
rect 525678 562170 525774 562226
rect 525154 562102 525774 562170
rect 525154 562046 525250 562102
rect 525306 562046 525374 562102
rect 525430 562046 525498 562102
rect 525554 562046 525622 562102
rect 525678 562046 525774 562102
rect 525154 561978 525774 562046
rect 525154 561922 525250 561978
rect 525306 561922 525374 561978
rect 525430 561922 525498 561978
rect 525554 561922 525622 561978
rect 525678 561922 525774 561978
rect 525154 544350 525774 561922
rect 525154 544294 525250 544350
rect 525306 544294 525374 544350
rect 525430 544294 525498 544350
rect 525554 544294 525622 544350
rect 525678 544294 525774 544350
rect 525154 544226 525774 544294
rect 525154 544170 525250 544226
rect 525306 544170 525374 544226
rect 525430 544170 525498 544226
rect 525554 544170 525622 544226
rect 525678 544170 525774 544226
rect 525154 544102 525774 544170
rect 525154 544046 525250 544102
rect 525306 544046 525374 544102
rect 525430 544046 525498 544102
rect 525554 544046 525622 544102
rect 525678 544046 525774 544102
rect 525154 543978 525774 544046
rect 525154 543922 525250 543978
rect 525306 543922 525374 543978
rect 525430 543922 525498 543978
rect 525554 543922 525622 543978
rect 525678 543922 525774 543978
rect 525154 527750 525774 543922
rect 528874 598172 529494 598268
rect 528874 598116 528970 598172
rect 529026 598116 529094 598172
rect 529150 598116 529218 598172
rect 529274 598116 529342 598172
rect 529398 598116 529494 598172
rect 528874 598048 529494 598116
rect 528874 597992 528970 598048
rect 529026 597992 529094 598048
rect 529150 597992 529218 598048
rect 529274 597992 529342 598048
rect 529398 597992 529494 598048
rect 528874 597924 529494 597992
rect 528874 597868 528970 597924
rect 529026 597868 529094 597924
rect 529150 597868 529218 597924
rect 529274 597868 529342 597924
rect 529398 597868 529494 597924
rect 528874 597800 529494 597868
rect 528874 597744 528970 597800
rect 529026 597744 529094 597800
rect 529150 597744 529218 597800
rect 529274 597744 529342 597800
rect 529398 597744 529494 597800
rect 528874 586350 529494 597744
rect 528874 586294 528970 586350
rect 529026 586294 529094 586350
rect 529150 586294 529218 586350
rect 529274 586294 529342 586350
rect 529398 586294 529494 586350
rect 528874 586226 529494 586294
rect 528874 586170 528970 586226
rect 529026 586170 529094 586226
rect 529150 586170 529218 586226
rect 529274 586170 529342 586226
rect 529398 586170 529494 586226
rect 528874 586102 529494 586170
rect 528874 586046 528970 586102
rect 529026 586046 529094 586102
rect 529150 586046 529218 586102
rect 529274 586046 529342 586102
rect 529398 586046 529494 586102
rect 528874 585978 529494 586046
rect 528874 585922 528970 585978
rect 529026 585922 529094 585978
rect 529150 585922 529218 585978
rect 529274 585922 529342 585978
rect 529398 585922 529494 585978
rect 528874 568350 529494 585922
rect 528874 568294 528970 568350
rect 529026 568294 529094 568350
rect 529150 568294 529218 568350
rect 529274 568294 529342 568350
rect 529398 568294 529494 568350
rect 528874 568226 529494 568294
rect 528874 568170 528970 568226
rect 529026 568170 529094 568226
rect 529150 568170 529218 568226
rect 529274 568170 529342 568226
rect 529398 568170 529494 568226
rect 528874 568102 529494 568170
rect 528874 568046 528970 568102
rect 529026 568046 529094 568102
rect 529150 568046 529218 568102
rect 529274 568046 529342 568102
rect 529398 568046 529494 568102
rect 528874 567978 529494 568046
rect 528874 567922 528970 567978
rect 529026 567922 529094 567978
rect 529150 567922 529218 567978
rect 529274 567922 529342 567978
rect 529398 567922 529494 567978
rect 528874 550350 529494 567922
rect 528874 550294 528970 550350
rect 529026 550294 529094 550350
rect 529150 550294 529218 550350
rect 529274 550294 529342 550350
rect 529398 550294 529494 550350
rect 528874 550226 529494 550294
rect 528874 550170 528970 550226
rect 529026 550170 529094 550226
rect 529150 550170 529218 550226
rect 529274 550170 529342 550226
rect 529398 550170 529494 550226
rect 528874 550102 529494 550170
rect 528874 550046 528970 550102
rect 529026 550046 529094 550102
rect 529150 550046 529218 550102
rect 529274 550046 529342 550102
rect 529398 550046 529494 550102
rect 528874 549978 529494 550046
rect 528874 549922 528970 549978
rect 529026 549922 529094 549978
rect 529150 549922 529218 549978
rect 529274 549922 529342 549978
rect 529398 549922 529494 549978
rect 528874 532350 529494 549922
rect 528874 532294 528970 532350
rect 529026 532294 529094 532350
rect 529150 532294 529218 532350
rect 529274 532294 529342 532350
rect 529398 532294 529494 532350
rect 528874 532226 529494 532294
rect 528874 532170 528970 532226
rect 529026 532170 529094 532226
rect 529150 532170 529218 532226
rect 529274 532170 529342 532226
rect 529398 532170 529494 532226
rect 528874 532102 529494 532170
rect 528874 532046 528970 532102
rect 529026 532046 529094 532102
rect 529150 532046 529218 532102
rect 529274 532046 529342 532102
rect 529398 532046 529494 532102
rect 528874 531978 529494 532046
rect 528874 531922 528970 531978
rect 529026 531922 529094 531978
rect 529150 531922 529218 531978
rect 529274 531922 529342 531978
rect 529398 531922 529494 531978
rect 528874 527750 529494 531922
rect 543154 597212 543774 598268
rect 543154 597156 543250 597212
rect 543306 597156 543374 597212
rect 543430 597156 543498 597212
rect 543554 597156 543622 597212
rect 543678 597156 543774 597212
rect 543154 597088 543774 597156
rect 543154 597032 543250 597088
rect 543306 597032 543374 597088
rect 543430 597032 543498 597088
rect 543554 597032 543622 597088
rect 543678 597032 543774 597088
rect 543154 596964 543774 597032
rect 543154 596908 543250 596964
rect 543306 596908 543374 596964
rect 543430 596908 543498 596964
rect 543554 596908 543622 596964
rect 543678 596908 543774 596964
rect 543154 596840 543774 596908
rect 543154 596784 543250 596840
rect 543306 596784 543374 596840
rect 543430 596784 543498 596840
rect 543554 596784 543622 596840
rect 543678 596784 543774 596840
rect 543154 580350 543774 596784
rect 543154 580294 543250 580350
rect 543306 580294 543374 580350
rect 543430 580294 543498 580350
rect 543554 580294 543622 580350
rect 543678 580294 543774 580350
rect 543154 580226 543774 580294
rect 543154 580170 543250 580226
rect 543306 580170 543374 580226
rect 543430 580170 543498 580226
rect 543554 580170 543622 580226
rect 543678 580170 543774 580226
rect 543154 580102 543774 580170
rect 543154 580046 543250 580102
rect 543306 580046 543374 580102
rect 543430 580046 543498 580102
rect 543554 580046 543622 580102
rect 543678 580046 543774 580102
rect 543154 579978 543774 580046
rect 543154 579922 543250 579978
rect 543306 579922 543374 579978
rect 543430 579922 543498 579978
rect 543554 579922 543622 579978
rect 543678 579922 543774 579978
rect 543154 562350 543774 579922
rect 543154 562294 543250 562350
rect 543306 562294 543374 562350
rect 543430 562294 543498 562350
rect 543554 562294 543622 562350
rect 543678 562294 543774 562350
rect 543154 562226 543774 562294
rect 543154 562170 543250 562226
rect 543306 562170 543374 562226
rect 543430 562170 543498 562226
rect 543554 562170 543622 562226
rect 543678 562170 543774 562226
rect 543154 562102 543774 562170
rect 543154 562046 543250 562102
rect 543306 562046 543374 562102
rect 543430 562046 543498 562102
rect 543554 562046 543622 562102
rect 543678 562046 543774 562102
rect 543154 561978 543774 562046
rect 543154 561922 543250 561978
rect 543306 561922 543374 561978
rect 543430 561922 543498 561978
rect 543554 561922 543622 561978
rect 543678 561922 543774 561978
rect 543154 544350 543774 561922
rect 543154 544294 543250 544350
rect 543306 544294 543374 544350
rect 543430 544294 543498 544350
rect 543554 544294 543622 544350
rect 543678 544294 543774 544350
rect 543154 544226 543774 544294
rect 543154 544170 543250 544226
rect 543306 544170 543374 544226
rect 543430 544170 543498 544226
rect 543554 544170 543622 544226
rect 543678 544170 543774 544226
rect 543154 544102 543774 544170
rect 543154 544046 543250 544102
rect 543306 544046 543374 544102
rect 543430 544046 543498 544102
rect 543554 544046 543622 544102
rect 543678 544046 543774 544102
rect 543154 543978 543774 544046
rect 543154 543922 543250 543978
rect 543306 543922 543374 543978
rect 543430 543922 543498 543978
rect 543554 543922 543622 543978
rect 543678 543922 543774 543978
rect 543154 527750 543774 543922
rect 546874 598172 547494 598268
rect 546874 598116 546970 598172
rect 547026 598116 547094 598172
rect 547150 598116 547218 598172
rect 547274 598116 547342 598172
rect 547398 598116 547494 598172
rect 546874 598048 547494 598116
rect 546874 597992 546970 598048
rect 547026 597992 547094 598048
rect 547150 597992 547218 598048
rect 547274 597992 547342 598048
rect 547398 597992 547494 598048
rect 546874 597924 547494 597992
rect 546874 597868 546970 597924
rect 547026 597868 547094 597924
rect 547150 597868 547218 597924
rect 547274 597868 547342 597924
rect 547398 597868 547494 597924
rect 546874 597800 547494 597868
rect 546874 597744 546970 597800
rect 547026 597744 547094 597800
rect 547150 597744 547218 597800
rect 547274 597744 547342 597800
rect 547398 597744 547494 597800
rect 546874 586350 547494 597744
rect 546874 586294 546970 586350
rect 547026 586294 547094 586350
rect 547150 586294 547218 586350
rect 547274 586294 547342 586350
rect 547398 586294 547494 586350
rect 546874 586226 547494 586294
rect 546874 586170 546970 586226
rect 547026 586170 547094 586226
rect 547150 586170 547218 586226
rect 547274 586170 547342 586226
rect 547398 586170 547494 586226
rect 546874 586102 547494 586170
rect 546874 586046 546970 586102
rect 547026 586046 547094 586102
rect 547150 586046 547218 586102
rect 547274 586046 547342 586102
rect 547398 586046 547494 586102
rect 546874 585978 547494 586046
rect 546874 585922 546970 585978
rect 547026 585922 547094 585978
rect 547150 585922 547218 585978
rect 547274 585922 547342 585978
rect 547398 585922 547494 585978
rect 546874 568350 547494 585922
rect 546874 568294 546970 568350
rect 547026 568294 547094 568350
rect 547150 568294 547218 568350
rect 547274 568294 547342 568350
rect 547398 568294 547494 568350
rect 546874 568226 547494 568294
rect 546874 568170 546970 568226
rect 547026 568170 547094 568226
rect 547150 568170 547218 568226
rect 547274 568170 547342 568226
rect 547398 568170 547494 568226
rect 546874 568102 547494 568170
rect 546874 568046 546970 568102
rect 547026 568046 547094 568102
rect 547150 568046 547218 568102
rect 547274 568046 547342 568102
rect 547398 568046 547494 568102
rect 546874 567978 547494 568046
rect 546874 567922 546970 567978
rect 547026 567922 547094 567978
rect 547150 567922 547218 567978
rect 547274 567922 547342 567978
rect 547398 567922 547494 567978
rect 546874 550350 547494 567922
rect 546874 550294 546970 550350
rect 547026 550294 547094 550350
rect 547150 550294 547218 550350
rect 547274 550294 547342 550350
rect 547398 550294 547494 550350
rect 546874 550226 547494 550294
rect 546874 550170 546970 550226
rect 547026 550170 547094 550226
rect 547150 550170 547218 550226
rect 547274 550170 547342 550226
rect 547398 550170 547494 550226
rect 546874 550102 547494 550170
rect 546874 550046 546970 550102
rect 547026 550046 547094 550102
rect 547150 550046 547218 550102
rect 547274 550046 547342 550102
rect 547398 550046 547494 550102
rect 546874 549978 547494 550046
rect 546874 549922 546970 549978
rect 547026 549922 547094 549978
rect 547150 549922 547218 549978
rect 547274 549922 547342 549978
rect 547398 549922 547494 549978
rect 546874 532350 547494 549922
rect 546874 532294 546970 532350
rect 547026 532294 547094 532350
rect 547150 532294 547218 532350
rect 547274 532294 547342 532350
rect 547398 532294 547494 532350
rect 546874 532226 547494 532294
rect 546874 532170 546970 532226
rect 547026 532170 547094 532226
rect 547150 532170 547218 532226
rect 547274 532170 547342 532226
rect 547398 532170 547494 532226
rect 546874 532102 547494 532170
rect 546874 532046 546970 532102
rect 547026 532046 547094 532102
rect 547150 532046 547218 532102
rect 547274 532046 547342 532102
rect 547398 532046 547494 532102
rect 546874 531978 547494 532046
rect 546874 531922 546970 531978
rect 547026 531922 547094 531978
rect 547150 531922 547218 531978
rect 547274 531922 547342 531978
rect 547398 531922 547494 531978
rect 546874 527750 547494 531922
rect 561154 597212 561774 598268
rect 561154 597156 561250 597212
rect 561306 597156 561374 597212
rect 561430 597156 561498 597212
rect 561554 597156 561622 597212
rect 561678 597156 561774 597212
rect 561154 597088 561774 597156
rect 561154 597032 561250 597088
rect 561306 597032 561374 597088
rect 561430 597032 561498 597088
rect 561554 597032 561622 597088
rect 561678 597032 561774 597088
rect 561154 596964 561774 597032
rect 561154 596908 561250 596964
rect 561306 596908 561374 596964
rect 561430 596908 561498 596964
rect 561554 596908 561622 596964
rect 561678 596908 561774 596964
rect 561154 596840 561774 596908
rect 561154 596784 561250 596840
rect 561306 596784 561374 596840
rect 561430 596784 561498 596840
rect 561554 596784 561622 596840
rect 561678 596784 561774 596840
rect 561154 580350 561774 596784
rect 561154 580294 561250 580350
rect 561306 580294 561374 580350
rect 561430 580294 561498 580350
rect 561554 580294 561622 580350
rect 561678 580294 561774 580350
rect 561154 580226 561774 580294
rect 561154 580170 561250 580226
rect 561306 580170 561374 580226
rect 561430 580170 561498 580226
rect 561554 580170 561622 580226
rect 561678 580170 561774 580226
rect 561154 580102 561774 580170
rect 561154 580046 561250 580102
rect 561306 580046 561374 580102
rect 561430 580046 561498 580102
rect 561554 580046 561622 580102
rect 561678 580046 561774 580102
rect 561154 579978 561774 580046
rect 561154 579922 561250 579978
rect 561306 579922 561374 579978
rect 561430 579922 561498 579978
rect 561554 579922 561622 579978
rect 561678 579922 561774 579978
rect 561154 562350 561774 579922
rect 561154 562294 561250 562350
rect 561306 562294 561374 562350
rect 561430 562294 561498 562350
rect 561554 562294 561622 562350
rect 561678 562294 561774 562350
rect 561154 562226 561774 562294
rect 561154 562170 561250 562226
rect 561306 562170 561374 562226
rect 561430 562170 561498 562226
rect 561554 562170 561622 562226
rect 561678 562170 561774 562226
rect 561154 562102 561774 562170
rect 561154 562046 561250 562102
rect 561306 562046 561374 562102
rect 561430 562046 561498 562102
rect 561554 562046 561622 562102
rect 561678 562046 561774 562102
rect 561154 561978 561774 562046
rect 561154 561922 561250 561978
rect 561306 561922 561374 561978
rect 561430 561922 561498 561978
rect 561554 561922 561622 561978
rect 561678 561922 561774 561978
rect 561154 544350 561774 561922
rect 561154 544294 561250 544350
rect 561306 544294 561374 544350
rect 561430 544294 561498 544350
rect 561554 544294 561622 544350
rect 561678 544294 561774 544350
rect 561154 544226 561774 544294
rect 561154 544170 561250 544226
rect 561306 544170 561374 544226
rect 561430 544170 561498 544226
rect 561554 544170 561622 544226
rect 561678 544170 561774 544226
rect 561154 544102 561774 544170
rect 561154 544046 561250 544102
rect 561306 544046 561374 544102
rect 561430 544046 561498 544102
rect 561554 544046 561622 544102
rect 561678 544046 561774 544102
rect 561154 543978 561774 544046
rect 561154 543922 561250 543978
rect 561306 543922 561374 543978
rect 561430 543922 561498 543978
rect 561554 543922 561622 543978
rect 561678 543922 561774 543978
rect 111154 526294 111250 526350
rect 111306 526294 111374 526350
rect 111430 526294 111498 526350
rect 111554 526294 111622 526350
rect 111678 526294 111774 526350
rect 561154 526350 561774 543922
rect 111154 526226 111774 526294
rect 111154 526170 111250 526226
rect 111306 526170 111374 526226
rect 111430 526170 111498 526226
rect 111554 526170 111622 526226
rect 111678 526170 111774 526226
rect 111154 526102 111774 526170
rect 111154 526046 111250 526102
rect 111306 526046 111374 526102
rect 111430 526046 111498 526102
rect 111554 526046 111622 526102
rect 111678 526046 111774 526102
rect 111154 525978 111774 526046
rect 111154 525922 111250 525978
rect 111306 525922 111374 525978
rect 111430 525922 111498 525978
rect 111554 525922 111622 525978
rect 111678 525922 111774 525978
rect 96874 514294 96970 514350
rect 97026 514294 97094 514350
rect 97150 514294 97218 514350
rect 97274 514294 97342 514350
rect 97398 514294 97494 514350
rect 96874 514226 97494 514294
rect 96874 514170 96970 514226
rect 97026 514170 97094 514226
rect 97150 514170 97218 514226
rect 97274 514170 97342 514226
rect 97398 514170 97494 514226
rect 96874 514102 97494 514170
rect 96874 514046 96970 514102
rect 97026 514046 97094 514102
rect 97150 514046 97218 514102
rect 97274 514046 97342 514102
rect 97398 514046 97494 514102
rect 96874 513978 97494 514046
rect 96874 513922 96970 513978
rect 97026 513922 97094 513978
rect 97150 513922 97218 513978
rect 97274 513922 97342 513978
rect 97398 513922 97494 513978
rect 96874 496350 97494 513922
rect 100528 514350 100848 514384
rect 100528 514294 100598 514350
rect 100654 514294 100722 514350
rect 100778 514294 100848 514350
rect 100528 514226 100848 514294
rect 100528 514170 100598 514226
rect 100654 514170 100722 514226
rect 100778 514170 100848 514226
rect 100528 514102 100848 514170
rect 100528 514046 100598 514102
rect 100654 514046 100722 514102
rect 100778 514046 100848 514102
rect 100528 513978 100848 514046
rect 100528 513922 100598 513978
rect 100654 513922 100722 513978
rect 100778 513922 100848 513978
rect 100528 513888 100848 513922
rect 111154 508350 111774 525922
rect 115888 526293 116208 526332
rect 115888 526237 115958 526293
rect 116014 526237 116082 526293
rect 116138 526237 116208 526293
rect 115888 526169 116208 526237
rect 115888 526113 115958 526169
rect 116014 526113 116082 526169
rect 116138 526113 116208 526169
rect 115888 526045 116208 526113
rect 115888 525989 115958 526045
rect 116014 525989 116082 526045
rect 116138 525989 116208 526045
rect 115888 525921 116208 525989
rect 115888 525865 115958 525921
rect 116014 525865 116082 525921
rect 116138 525865 116208 525921
rect 115888 525826 116208 525865
rect 146608 526293 146928 526332
rect 146608 526237 146678 526293
rect 146734 526237 146802 526293
rect 146858 526237 146928 526293
rect 146608 526169 146928 526237
rect 146608 526113 146678 526169
rect 146734 526113 146802 526169
rect 146858 526113 146928 526169
rect 146608 526045 146928 526113
rect 146608 525989 146678 526045
rect 146734 525989 146802 526045
rect 146858 525989 146928 526045
rect 146608 525921 146928 525989
rect 146608 525865 146678 525921
rect 146734 525865 146802 525921
rect 146858 525865 146928 525921
rect 146608 525826 146928 525865
rect 177328 526293 177648 526332
rect 177328 526237 177398 526293
rect 177454 526237 177522 526293
rect 177578 526237 177648 526293
rect 177328 526169 177648 526237
rect 177328 526113 177398 526169
rect 177454 526113 177522 526169
rect 177578 526113 177648 526169
rect 177328 526045 177648 526113
rect 177328 525989 177398 526045
rect 177454 525989 177522 526045
rect 177578 525989 177648 526045
rect 177328 525921 177648 525989
rect 177328 525865 177398 525921
rect 177454 525865 177522 525921
rect 177578 525865 177648 525921
rect 177328 525826 177648 525865
rect 208048 526293 208368 526332
rect 208048 526237 208118 526293
rect 208174 526237 208242 526293
rect 208298 526237 208368 526293
rect 208048 526169 208368 526237
rect 208048 526113 208118 526169
rect 208174 526113 208242 526169
rect 208298 526113 208368 526169
rect 208048 526045 208368 526113
rect 208048 525989 208118 526045
rect 208174 525989 208242 526045
rect 208298 525989 208368 526045
rect 208048 525921 208368 525989
rect 208048 525865 208118 525921
rect 208174 525865 208242 525921
rect 208298 525865 208368 525921
rect 208048 525826 208368 525865
rect 238768 526293 239088 526332
rect 238768 526237 238838 526293
rect 238894 526237 238962 526293
rect 239018 526237 239088 526293
rect 238768 526169 239088 526237
rect 238768 526113 238838 526169
rect 238894 526113 238962 526169
rect 239018 526113 239088 526169
rect 238768 526045 239088 526113
rect 238768 525989 238838 526045
rect 238894 525989 238962 526045
rect 239018 525989 239088 526045
rect 238768 525921 239088 525989
rect 238768 525865 238838 525921
rect 238894 525865 238962 525921
rect 239018 525865 239088 525921
rect 238768 525826 239088 525865
rect 269488 526293 269808 526332
rect 269488 526237 269558 526293
rect 269614 526237 269682 526293
rect 269738 526237 269808 526293
rect 269488 526169 269808 526237
rect 269488 526113 269558 526169
rect 269614 526113 269682 526169
rect 269738 526113 269808 526169
rect 269488 526045 269808 526113
rect 269488 525989 269558 526045
rect 269614 525989 269682 526045
rect 269738 525989 269808 526045
rect 269488 525921 269808 525989
rect 269488 525865 269558 525921
rect 269614 525865 269682 525921
rect 269738 525865 269808 525921
rect 269488 525826 269808 525865
rect 300208 526293 300528 526332
rect 300208 526237 300278 526293
rect 300334 526237 300402 526293
rect 300458 526237 300528 526293
rect 300208 526169 300528 526237
rect 300208 526113 300278 526169
rect 300334 526113 300402 526169
rect 300458 526113 300528 526169
rect 300208 526045 300528 526113
rect 300208 525989 300278 526045
rect 300334 525989 300402 526045
rect 300458 525989 300528 526045
rect 300208 525921 300528 525989
rect 300208 525865 300278 525921
rect 300334 525865 300402 525921
rect 300458 525865 300528 525921
rect 300208 525826 300528 525865
rect 330928 526293 331248 526332
rect 330928 526237 330998 526293
rect 331054 526237 331122 526293
rect 331178 526237 331248 526293
rect 330928 526169 331248 526237
rect 330928 526113 330998 526169
rect 331054 526113 331122 526169
rect 331178 526113 331248 526169
rect 330928 526045 331248 526113
rect 330928 525989 330998 526045
rect 331054 525989 331122 526045
rect 331178 525989 331248 526045
rect 330928 525921 331248 525989
rect 330928 525865 330998 525921
rect 331054 525865 331122 525921
rect 331178 525865 331248 525921
rect 330928 525826 331248 525865
rect 361648 526293 361968 526332
rect 361648 526237 361718 526293
rect 361774 526237 361842 526293
rect 361898 526237 361968 526293
rect 361648 526169 361968 526237
rect 361648 526113 361718 526169
rect 361774 526113 361842 526169
rect 361898 526113 361968 526169
rect 361648 526045 361968 526113
rect 361648 525989 361718 526045
rect 361774 525989 361842 526045
rect 361898 525989 361968 526045
rect 361648 525921 361968 525989
rect 361648 525865 361718 525921
rect 361774 525865 361842 525921
rect 361898 525865 361968 525921
rect 361648 525826 361968 525865
rect 392368 526293 392688 526332
rect 392368 526237 392438 526293
rect 392494 526237 392562 526293
rect 392618 526237 392688 526293
rect 392368 526169 392688 526237
rect 392368 526113 392438 526169
rect 392494 526113 392562 526169
rect 392618 526113 392688 526169
rect 392368 526045 392688 526113
rect 392368 525989 392438 526045
rect 392494 525989 392562 526045
rect 392618 525989 392688 526045
rect 392368 525921 392688 525989
rect 392368 525865 392438 525921
rect 392494 525865 392562 525921
rect 392618 525865 392688 525921
rect 392368 525826 392688 525865
rect 423088 526293 423408 526332
rect 423088 526237 423158 526293
rect 423214 526237 423282 526293
rect 423338 526237 423408 526293
rect 423088 526169 423408 526237
rect 423088 526113 423158 526169
rect 423214 526113 423282 526169
rect 423338 526113 423408 526169
rect 423088 526045 423408 526113
rect 423088 525989 423158 526045
rect 423214 525989 423282 526045
rect 423338 525989 423408 526045
rect 423088 525921 423408 525989
rect 423088 525865 423158 525921
rect 423214 525865 423282 525921
rect 423338 525865 423408 525921
rect 423088 525826 423408 525865
rect 453808 526293 454128 526332
rect 453808 526237 453878 526293
rect 453934 526237 454002 526293
rect 454058 526237 454128 526293
rect 453808 526169 454128 526237
rect 453808 526113 453878 526169
rect 453934 526113 454002 526169
rect 454058 526113 454128 526169
rect 453808 526045 454128 526113
rect 453808 525989 453878 526045
rect 453934 525989 454002 526045
rect 454058 525989 454128 526045
rect 453808 525921 454128 525989
rect 453808 525865 453878 525921
rect 453934 525865 454002 525921
rect 454058 525865 454128 525921
rect 453808 525826 454128 525865
rect 484528 526293 484848 526332
rect 484528 526237 484598 526293
rect 484654 526237 484722 526293
rect 484778 526237 484848 526293
rect 484528 526169 484848 526237
rect 484528 526113 484598 526169
rect 484654 526113 484722 526169
rect 484778 526113 484848 526169
rect 484528 526045 484848 526113
rect 484528 525989 484598 526045
rect 484654 525989 484722 526045
rect 484778 525989 484848 526045
rect 484528 525921 484848 525989
rect 484528 525865 484598 525921
rect 484654 525865 484722 525921
rect 484778 525865 484848 525921
rect 484528 525826 484848 525865
rect 515248 526293 515568 526332
rect 515248 526237 515318 526293
rect 515374 526237 515442 526293
rect 515498 526237 515568 526293
rect 515248 526169 515568 526237
rect 515248 526113 515318 526169
rect 515374 526113 515442 526169
rect 515498 526113 515568 526169
rect 515248 526045 515568 526113
rect 515248 525989 515318 526045
rect 515374 525989 515442 526045
rect 515498 525989 515568 526045
rect 515248 525921 515568 525989
rect 515248 525865 515318 525921
rect 515374 525865 515442 525921
rect 515498 525865 515568 525921
rect 515248 525826 515568 525865
rect 545968 526293 546288 526332
rect 545968 526237 546038 526293
rect 546094 526237 546162 526293
rect 546218 526237 546288 526293
rect 545968 526169 546288 526237
rect 545968 526113 546038 526169
rect 546094 526113 546162 526169
rect 546218 526113 546288 526169
rect 545968 526045 546288 526113
rect 545968 525989 546038 526045
rect 546094 525989 546162 526045
rect 546218 525989 546288 526045
rect 545968 525921 546288 525989
rect 545968 525865 546038 525921
rect 546094 525865 546162 525921
rect 546218 525865 546288 525921
rect 545968 525826 546288 525865
rect 561154 526294 561250 526350
rect 561306 526294 561374 526350
rect 561430 526294 561498 526350
rect 561554 526294 561622 526350
rect 561678 526294 561774 526350
rect 561154 526226 561774 526294
rect 561154 526170 561250 526226
rect 561306 526170 561374 526226
rect 561430 526170 561498 526226
rect 561554 526170 561622 526226
rect 561678 526170 561774 526226
rect 561154 526102 561774 526170
rect 561154 526046 561250 526102
rect 561306 526046 561374 526102
rect 561430 526046 561498 526102
rect 561554 526046 561622 526102
rect 561678 526046 561774 526102
rect 561154 525978 561774 526046
rect 561154 525922 561250 525978
rect 561306 525922 561374 525978
rect 561430 525922 561498 525978
rect 561554 525922 561622 525978
rect 561678 525922 561774 525978
rect 131248 514350 131568 514384
rect 131248 514294 131318 514350
rect 131374 514294 131442 514350
rect 131498 514294 131568 514350
rect 131248 514226 131568 514294
rect 131248 514170 131318 514226
rect 131374 514170 131442 514226
rect 131498 514170 131568 514226
rect 131248 514102 131568 514170
rect 131248 514046 131318 514102
rect 131374 514046 131442 514102
rect 131498 514046 131568 514102
rect 131248 513978 131568 514046
rect 131248 513922 131318 513978
rect 131374 513922 131442 513978
rect 131498 513922 131568 513978
rect 131248 513888 131568 513922
rect 161968 514350 162288 514384
rect 161968 514294 162038 514350
rect 162094 514294 162162 514350
rect 162218 514294 162288 514350
rect 161968 514226 162288 514294
rect 161968 514170 162038 514226
rect 162094 514170 162162 514226
rect 162218 514170 162288 514226
rect 161968 514102 162288 514170
rect 161968 514046 162038 514102
rect 162094 514046 162162 514102
rect 162218 514046 162288 514102
rect 161968 513978 162288 514046
rect 161968 513922 162038 513978
rect 162094 513922 162162 513978
rect 162218 513922 162288 513978
rect 161968 513888 162288 513922
rect 192688 514350 193008 514384
rect 192688 514294 192758 514350
rect 192814 514294 192882 514350
rect 192938 514294 193008 514350
rect 192688 514226 193008 514294
rect 192688 514170 192758 514226
rect 192814 514170 192882 514226
rect 192938 514170 193008 514226
rect 192688 514102 193008 514170
rect 192688 514046 192758 514102
rect 192814 514046 192882 514102
rect 192938 514046 193008 514102
rect 192688 513978 193008 514046
rect 192688 513922 192758 513978
rect 192814 513922 192882 513978
rect 192938 513922 193008 513978
rect 192688 513888 193008 513922
rect 223408 514350 223728 514384
rect 223408 514294 223478 514350
rect 223534 514294 223602 514350
rect 223658 514294 223728 514350
rect 223408 514226 223728 514294
rect 223408 514170 223478 514226
rect 223534 514170 223602 514226
rect 223658 514170 223728 514226
rect 223408 514102 223728 514170
rect 223408 514046 223478 514102
rect 223534 514046 223602 514102
rect 223658 514046 223728 514102
rect 223408 513978 223728 514046
rect 223408 513922 223478 513978
rect 223534 513922 223602 513978
rect 223658 513922 223728 513978
rect 223408 513888 223728 513922
rect 254128 514350 254448 514384
rect 254128 514294 254198 514350
rect 254254 514294 254322 514350
rect 254378 514294 254448 514350
rect 254128 514226 254448 514294
rect 254128 514170 254198 514226
rect 254254 514170 254322 514226
rect 254378 514170 254448 514226
rect 254128 514102 254448 514170
rect 254128 514046 254198 514102
rect 254254 514046 254322 514102
rect 254378 514046 254448 514102
rect 254128 513978 254448 514046
rect 254128 513922 254198 513978
rect 254254 513922 254322 513978
rect 254378 513922 254448 513978
rect 254128 513888 254448 513922
rect 284848 514350 285168 514384
rect 284848 514294 284918 514350
rect 284974 514294 285042 514350
rect 285098 514294 285168 514350
rect 284848 514226 285168 514294
rect 284848 514170 284918 514226
rect 284974 514170 285042 514226
rect 285098 514170 285168 514226
rect 284848 514102 285168 514170
rect 284848 514046 284918 514102
rect 284974 514046 285042 514102
rect 285098 514046 285168 514102
rect 284848 513978 285168 514046
rect 284848 513922 284918 513978
rect 284974 513922 285042 513978
rect 285098 513922 285168 513978
rect 284848 513888 285168 513922
rect 315568 514350 315888 514384
rect 315568 514294 315638 514350
rect 315694 514294 315762 514350
rect 315818 514294 315888 514350
rect 315568 514226 315888 514294
rect 315568 514170 315638 514226
rect 315694 514170 315762 514226
rect 315818 514170 315888 514226
rect 315568 514102 315888 514170
rect 315568 514046 315638 514102
rect 315694 514046 315762 514102
rect 315818 514046 315888 514102
rect 315568 513978 315888 514046
rect 315568 513922 315638 513978
rect 315694 513922 315762 513978
rect 315818 513922 315888 513978
rect 315568 513888 315888 513922
rect 346288 514350 346608 514384
rect 346288 514294 346358 514350
rect 346414 514294 346482 514350
rect 346538 514294 346608 514350
rect 346288 514226 346608 514294
rect 346288 514170 346358 514226
rect 346414 514170 346482 514226
rect 346538 514170 346608 514226
rect 346288 514102 346608 514170
rect 346288 514046 346358 514102
rect 346414 514046 346482 514102
rect 346538 514046 346608 514102
rect 346288 513978 346608 514046
rect 346288 513922 346358 513978
rect 346414 513922 346482 513978
rect 346538 513922 346608 513978
rect 346288 513888 346608 513922
rect 377008 514350 377328 514384
rect 377008 514294 377078 514350
rect 377134 514294 377202 514350
rect 377258 514294 377328 514350
rect 377008 514226 377328 514294
rect 377008 514170 377078 514226
rect 377134 514170 377202 514226
rect 377258 514170 377328 514226
rect 377008 514102 377328 514170
rect 377008 514046 377078 514102
rect 377134 514046 377202 514102
rect 377258 514046 377328 514102
rect 377008 513978 377328 514046
rect 377008 513922 377078 513978
rect 377134 513922 377202 513978
rect 377258 513922 377328 513978
rect 377008 513888 377328 513922
rect 407728 514350 408048 514384
rect 407728 514294 407798 514350
rect 407854 514294 407922 514350
rect 407978 514294 408048 514350
rect 407728 514226 408048 514294
rect 407728 514170 407798 514226
rect 407854 514170 407922 514226
rect 407978 514170 408048 514226
rect 407728 514102 408048 514170
rect 407728 514046 407798 514102
rect 407854 514046 407922 514102
rect 407978 514046 408048 514102
rect 407728 513978 408048 514046
rect 407728 513922 407798 513978
rect 407854 513922 407922 513978
rect 407978 513922 408048 513978
rect 407728 513888 408048 513922
rect 438448 514350 438768 514384
rect 438448 514294 438518 514350
rect 438574 514294 438642 514350
rect 438698 514294 438768 514350
rect 438448 514226 438768 514294
rect 438448 514170 438518 514226
rect 438574 514170 438642 514226
rect 438698 514170 438768 514226
rect 438448 514102 438768 514170
rect 438448 514046 438518 514102
rect 438574 514046 438642 514102
rect 438698 514046 438768 514102
rect 438448 513978 438768 514046
rect 438448 513922 438518 513978
rect 438574 513922 438642 513978
rect 438698 513922 438768 513978
rect 438448 513888 438768 513922
rect 469168 514350 469488 514384
rect 469168 514294 469238 514350
rect 469294 514294 469362 514350
rect 469418 514294 469488 514350
rect 469168 514226 469488 514294
rect 469168 514170 469238 514226
rect 469294 514170 469362 514226
rect 469418 514170 469488 514226
rect 469168 514102 469488 514170
rect 469168 514046 469238 514102
rect 469294 514046 469362 514102
rect 469418 514046 469488 514102
rect 469168 513978 469488 514046
rect 469168 513922 469238 513978
rect 469294 513922 469362 513978
rect 469418 513922 469488 513978
rect 469168 513888 469488 513922
rect 499888 514350 500208 514384
rect 499888 514294 499958 514350
rect 500014 514294 500082 514350
rect 500138 514294 500208 514350
rect 499888 514226 500208 514294
rect 499888 514170 499958 514226
rect 500014 514170 500082 514226
rect 500138 514170 500208 514226
rect 499888 514102 500208 514170
rect 499888 514046 499958 514102
rect 500014 514046 500082 514102
rect 500138 514046 500208 514102
rect 499888 513978 500208 514046
rect 499888 513922 499958 513978
rect 500014 513922 500082 513978
rect 500138 513922 500208 513978
rect 499888 513888 500208 513922
rect 530608 514350 530928 514384
rect 530608 514294 530678 514350
rect 530734 514294 530802 514350
rect 530858 514294 530928 514350
rect 530608 514226 530928 514294
rect 530608 514170 530678 514226
rect 530734 514170 530802 514226
rect 530858 514170 530928 514226
rect 530608 514102 530928 514170
rect 530608 514046 530678 514102
rect 530734 514046 530802 514102
rect 530858 514046 530928 514102
rect 530608 513978 530928 514046
rect 530608 513922 530678 513978
rect 530734 513922 530802 513978
rect 530858 513922 530928 513978
rect 530608 513888 530928 513922
rect 111154 508294 111250 508350
rect 111306 508294 111374 508350
rect 111430 508294 111498 508350
rect 111554 508294 111622 508350
rect 111678 508294 111774 508350
rect 111154 508226 111774 508294
rect 111154 508170 111250 508226
rect 111306 508170 111374 508226
rect 111430 508170 111498 508226
rect 111554 508170 111622 508226
rect 111678 508170 111774 508226
rect 111154 508102 111774 508170
rect 111154 508046 111250 508102
rect 111306 508046 111374 508102
rect 111430 508046 111498 508102
rect 111554 508046 111622 508102
rect 111678 508046 111774 508102
rect 111154 507978 111774 508046
rect 111154 507922 111250 507978
rect 111306 507922 111374 507978
rect 111430 507922 111498 507978
rect 111554 507922 111622 507978
rect 111678 507922 111774 507978
rect 96874 496294 96970 496350
rect 97026 496294 97094 496350
rect 97150 496294 97218 496350
rect 97274 496294 97342 496350
rect 97398 496294 97494 496350
rect 96874 496226 97494 496294
rect 96874 496170 96970 496226
rect 97026 496170 97094 496226
rect 97150 496170 97218 496226
rect 97274 496170 97342 496226
rect 97398 496170 97494 496226
rect 96874 496102 97494 496170
rect 96874 496046 96970 496102
rect 97026 496046 97094 496102
rect 97150 496046 97218 496102
rect 97274 496046 97342 496102
rect 97398 496046 97494 496102
rect 96874 495978 97494 496046
rect 96874 495922 96970 495978
rect 97026 495922 97094 495978
rect 97150 495922 97218 495978
rect 97274 495922 97342 495978
rect 97398 495922 97494 495978
rect 96874 478350 97494 495922
rect 100528 496350 100848 496384
rect 100528 496294 100598 496350
rect 100654 496294 100722 496350
rect 100778 496294 100848 496350
rect 100528 496226 100848 496294
rect 100528 496170 100598 496226
rect 100654 496170 100722 496226
rect 100778 496170 100848 496226
rect 100528 496102 100848 496170
rect 100528 496046 100598 496102
rect 100654 496046 100722 496102
rect 100778 496046 100848 496102
rect 100528 495978 100848 496046
rect 100528 495922 100598 495978
rect 100654 495922 100722 495978
rect 100778 495922 100848 495978
rect 100528 495888 100848 495922
rect 111154 490350 111774 507922
rect 115888 508350 116208 508384
rect 115888 508294 115958 508350
rect 116014 508294 116082 508350
rect 116138 508294 116208 508350
rect 115888 508226 116208 508294
rect 115888 508170 115958 508226
rect 116014 508170 116082 508226
rect 116138 508170 116208 508226
rect 115888 508102 116208 508170
rect 115888 508046 115958 508102
rect 116014 508046 116082 508102
rect 116138 508046 116208 508102
rect 115888 507978 116208 508046
rect 115888 507922 115958 507978
rect 116014 507922 116082 507978
rect 116138 507922 116208 507978
rect 115888 507888 116208 507922
rect 146608 508350 146928 508384
rect 146608 508294 146678 508350
rect 146734 508294 146802 508350
rect 146858 508294 146928 508350
rect 146608 508226 146928 508294
rect 146608 508170 146678 508226
rect 146734 508170 146802 508226
rect 146858 508170 146928 508226
rect 146608 508102 146928 508170
rect 146608 508046 146678 508102
rect 146734 508046 146802 508102
rect 146858 508046 146928 508102
rect 146608 507978 146928 508046
rect 146608 507922 146678 507978
rect 146734 507922 146802 507978
rect 146858 507922 146928 507978
rect 146608 507888 146928 507922
rect 177328 508350 177648 508384
rect 177328 508294 177398 508350
rect 177454 508294 177522 508350
rect 177578 508294 177648 508350
rect 177328 508226 177648 508294
rect 177328 508170 177398 508226
rect 177454 508170 177522 508226
rect 177578 508170 177648 508226
rect 177328 508102 177648 508170
rect 177328 508046 177398 508102
rect 177454 508046 177522 508102
rect 177578 508046 177648 508102
rect 177328 507978 177648 508046
rect 177328 507922 177398 507978
rect 177454 507922 177522 507978
rect 177578 507922 177648 507978
rect 177328 507888 177648 507922
rect 208048 508350 208368 508384
rect 208048 508294 208118 508350
rect 208174 508294 208242 508350
rect 208298 508294 208368 508350
rect 208048 508226 208368 508294
rect 208048 508170 208118 508226
rect 208174 508170 208242 508226
rect 208298 508170 208368 508226
rect 208048 508102 208368 508170
rect 208048 508046 208118 508102
rect 208174 508046 208242 508102
rect 208298 508046 208368 508102
rect 208048 507978 208368 508046
rect 208048 507922 208118 507978
rect 208174 507922 208242 507978
rect 208298 507922 208368 507978
rect 208048 507888 208368 507922
rect 238768 508350 239088 508384
rect 238768 508294 238838 508350
rect 238894 508294 238962 508350
rect 239018 508294 239088 508350
rect 238768 508226 239088 508294
rect 238768 508170 238838 508226
rect 238894 508170 238962 508226
rect 239018 508170 239088 508226
rect 238768 508102 239088 508170
rect 238768 508046 238838 508102
rect 238894 508046 238962 508102
rect 239018 508046 239088 508102
rect 238768 507978 239088 508046
rect 238768 507922 238838 507978
rect 238894 507922 238962 507978
rect 239018 507922 239088 507978
rect 238768 507888 239088 507922
rect 269488 508350 269808 508384
rect 269488 508294 269558 508350
rect 269614 508294 269682 508350
rect 269738 508294 269808 508350
rect 269488 508226 269808 508294
rect 269488 508170 269558 508226
rect 269614 508170 269682 508226
rect 269738 508170 269808 508226
rect 269488 508102 269808 508170
rect 269488 508046 269558 508102
rect 269614 508046 269682 508102
rect 269738 508046 269808 508102
rect 269488 507978 269808 508046
rect 269488 507922 269558 507978
rect 269614 507922 269682 507978
rect 269738 507922 269808 507978
rect 269488 507888 269808 507922
rect 300208 508350 300528 508384
rect 300208 508294 300278 508350
rect 300334 508294 300402 508350
rect 300458 508294 300528 508350
rect 300208 508226 300528 508294
rect 300208 508170 300278 508226
rect 300334 508170 300402 508226
rect 300458 508170 300528 508226
rect 300208 508102 300528 508170
rect 300208 508046 300278 508102
rect 300334 508046 300402 508102
rect 300458 508046 300528 508102
rect 300208 507978 300528 508046
rect 300208 507922 300278 507978
rect 300334 507922 300402 507978
rect 300458 507922 300528 507978
rect 300208 507888 300528 507922
rect 330928 508350 331248 508384
rect 330928 508294 330998 508350
rect 331054 508294 331122 508350
rect 331178 508294 331248 508350
rect 330928 508226 331248 508294
rect 330928 508170 330998 508226
rect 331054 508170 331122 508226
rect 331178 508170 331248 508226
rect 330928 508102 331248 508170
rect 330928 508046 330998 508102
rect 331054 508046 331122 508102
rect 331178 508046 331248 508102
rect 330928 507978 331248 508046
rect 330928 507922 330998 507978
rect 331054 507922 331122 507978
rect 331178 507922 331248 507978
rect 330928 507888 331248 507922
rect 361648 508350 361968 508384
rect 361648 508294 361718 508350
rect 361774 508294 361842 508350
rect 361898 508294 361968 508350
rect 361648 508226 361968 508294
rect 361648 508170 361718 508226
rect 361774 508170 361842 508226
rect 361898 508170 361968 508226
rect 361648 508102 361968 508170
rect 361648 508046 361718 508102
rect 361774 508046 361842 508102
rect 361898 508046 361968 508102
rect 361648 507978 361968 508046
rect 361648 507922 361718 507978
rect 361774 507922 361842 507978
rect 361898 507922 361968 507978
rect 361648 507888 361968 507922
rect 392368 508350 392688 508384
rect 392368 508294 392438 508350
rect 392494 508294 392562 508350
rect 392618 508294 392688 508350
rect 392368 508226 392688 508294
rect 392368 508170 392438 508226
rect 392494 508170 392562 508226
rect 392618 508170 392688 508226
rect 392368 508102 392688 508170
rect 392368 508046 392438 508102
rect 392494 508046 392562 508102
rect 392618 508046 392688 508102
rect 392368 507978 392688 508046
rect 392368 507922 392438 507978
rect 392494 507922 392562 507978
rect 392618 507922 392688 507978
rect 392368 507888 392688 507922
rect 423088 508350 423408 508384
rect 423088 508294 423158 508350
rect 423214 508294 423282 508350
rect 423338 508294 423408 508350
rect 423088 508226 423408 508294
rect 423088 508170 423158 508226
rect 423214 508170 423282 508226
rect 423338 508170 423408 508226
rect 423088 508102 423408 508170
rect 423088 508046 423158 508102
rect 423214 508046 423282 508102
rect 423338 508046 423408 508102
rect 423088 507978 423408 508046
rect 423088 507922 423158 507978
rect 423214 507922 423282 507978
rect 423338 507922 423408 507978
rect 423088 507888 423408 507922
rect 453808 508350 454128 508384
rect 453808 508294 453878 508350
rect 453934 508294 454002 508350
rect 454058 508294 454128 508350
rect 453808 508226 454128 508294
rect 453808 508170 453878 508226
rect 453934 508170 454002 508226
rect 454058 508170 454128 508226
rect 453808 508102 454128 508170
rect 453808 508046 453878 508102
rect 453934 508046 454002 508102
rect 454058 508046 454128 508102
rect 453808 507978 454128 508046
rect 453808 507922 453878 507978
rect 453934 507922 454002 507978
rect 454058 507922 454128 507978
rect 453808 507888 454128 507922
rect 484528 508350 484848 508384
rect 484528 508294 484598 508350
rect 484654 508294 484722 508350
rect 484778 508294 484848 508350
rect 484528 508226 484848 508294
rect 484528 508170 484598 508226
rect 484654 508170 484722 508226
rect 484778 508170 484848 508226
rect 484528 508102 484848 508170
rect 484528 508046 484598 508102
rect 484654 508046 484722 508102
rect 484778 508046 484848 508102
rect 484528 507978 484848 508046
rect 484528 507922 484598 507978
rect 484654 507922 484722 507978
rect 484778 507922 484848 507978
rect 484528 507888 484848 507922
rect 515248 508350 515568 508384
rect 515248 508294 515318 508350
rect 515374 508294 515442 508350
rect 515498 508294 515568 508350
rect 515248 508226 515568 508294
rect 515248 508170 515318 508226
rect 515374 508170 515442 508226
rect 515498 508170 515568 508226
rect 515248 508102 515568 508170
rect 515248 508046 515318 508102
rect 515374 508046 515442 508102
rect 515498 508046 515568 508102
rect 515248 507978 515568 508046
rect 515248 507922 515318 507978
rect 515374 507922 515442 507978
rect 515498 507922 515568 507978
rect 515248 507888 515568 507922
rect 545968 508350 546288 508384
rect 545968 508294 546038 508350
rect 546094 508294 546162 508350
rect 546218 508294 546288 508350
rect 545968 508226 546288 508294
rect 545968 508170 546038 508226
rect 546094 508170 546162 508226
rect 546218 508170 546288 508226
rect 545968 508102 546288 508170
rect 545968 508046 546038 508102
rect 546094 508046 546162 508102
rect 546218 508046 546288 508102
rect 545968 507978 546288 508046
rect 545968 507922 546038 507978
rect 546094 507922 546162 507978
rect 546218 507922 546288 507978
rect 545968 507888 546288 507922
rect 561154 508350 561774 525922
rect 561154 508294 561250 508350
rect 561306 508294 561374 508350
rect 561430 508294 561498 508350
rect 561554 508294 561622 508350
rect 561678 508294 561774 508350
rect 561154 508226 561774 508294
rect 561154 508170 561250 508226
rect 561306 508170 561374 508226
rect 561430 508170 561498 508226
rect 561554 508170 561622 508226
rect 561678 508170 561774 508226
rect 561154 508102 561774 508170
rect 561154 508046 561250 508102
rect 561306 508046 561374 508102
rect 561430 508046 561498 508102
rect 561554 508046 561622 508102
rect 561678 508046 561774 508102
rect 561154 507978 561774 508046
rect 561154 507922 561250 507978
rect 561306 507922 561374 507978
rect 561430 507922 561498 507978
rect 561554 507922 561622 507978
rect 561678 507922 561774 507978
rect 131248 496350 131568 496384
rect 131248 496294 131318 496350
rect 131374 496294 131442 496350
rect 131498 496294 131568 496350
rect 131248 496226 131568 496294
rect 131248 496170 131318 496226
rect 131374 496170 131442 496226
rect 131498 496170 131568 496226
rect 131248 496102 131568 496170
rect 131248 496046 131318 496102
rect 131374 496046 131442 496102
rect 131498 496046 131568 496102
rect 131248 495978 131568 496046
rect 131248 495922 131318 495978
rect 131374 495922 131442 495978
rect 131498 495922 131568 495978
rect 131248 495888 131568 495922
rect 161968 496350 162288 496384
rect 161968 496294 162038 496350
rect 162094 496294 162162 496350
rect 162218 496294 162288 496350
rect 161968 496226 162288 496294
rect 161968 496170 162038 496226
rect 162094 496170 162162 496226
rect 162218 496170 162288 496226
rect 161968 496102 162288 496170
rect 161968 496046 162038 496102
rect 162094 496046 162162 496102
rect 162218 496046 162288 496102
rect 161968 495978 162288 496046
rect 161968 495922 162038 495978
rect 162094 495922 162162 495978
rect 162218 495922 162288 495978
rect 161968 495888 162288 495922
rect 192688 496350 193008 496384
rect 192688 496294 192758 496350
rect 192814 496294 192882 496350
rect 192938 496294 193008 496350
rect 192688 496226 193008 496294
rect 192688 496170 192758 496226
rect 192814 496170 192882 496226
rect 192938 496170 193008 496226
rect 192688 496102 193008 496170
rect 192688 496046 192758 496102
rect 192814 496046 192882 496102
rect 192938 496046 193008 496102
rect 192688 495978 193008 496046
rect 192688 495922 192758 495978
rect 192814 495922 192882 495978
rect 192938 495922 193008 495978
rect 192688 495888 193008 495922
rect 223408 496350 223728 496384
rect 223408 496294 223478 496350
rect 223534 496294 223602 496350
rect 223658 496294 223728 496350
rect 223408 496226 223728 496294
rect 223408 496170 223478 496226
rect 223534 496170 223602 496226
rect 223658 496170 223728 496226
rect 223408 496102 223728 496170
rect 223408 496046 223478 496102
rect 223534 496046 223602 496102
rect 223658 496046 223728 496102
rect 223408 495978 223728 496046
rect 223408 495922 223478 495978
rect 223534 495922 223602 495978
rect 223658 495922 223728 495978
rect 223408 495888 223728 495922
rect 254128 496350 254448 496384
rect 254128 496294 254198 496350
rect 254254 496294 254322 496350
rect 254378 496294 254448 496350
rect 254128 496226 254448 496294
rect 254128 496170 254198 496226
rect 254254 496170 254322 496226
rect 254378 496170 254448 496226
rect 254128 496102 254448 496170
rect 254128 496046 254198 496102
rect 254254 496046 254322 496102
rect 254378 496046 254448 496102
rect 254128 495978 254448 496046
rect 254128 495922 254198 495978
rect 254254 495922 254322 495978
rect 254378 495922 254448 495978
rect 254128 495888 254448 495922
rect 284848 496350 285168 496384
rect 284848 496294 284918 496350
rect 284974 496294 285042 496350
rect 285098 496294 285168 496350
rect 284848 496226 285168 496294
rect 284848 496170 284918 496226
rect 284974 496170 285042 496226
rect 285098 496170 285168 496226
rect 284848 496102 285168 496170
rect 284848 496046 284918 496102
rect 284974 496046 285042 496102
rect 285098 496046 285168 496102
rect 284848 495978 285168 496046
rect 284848 495922 284918 495978
rect 284974 495922 285042 495978
rect 285098 495922 285168 495978
rect 284848 495888 285168 495922
rect 315568 496350 315888 496384
rect 315568 496294 315638 496350
rect 315694 496294 315762 496350
rect 315818 496294 315888 496350
rect 315568 496226 315888 496294
rect 315568 496170 315638 496226
rect 315694 496170 315762 496226
rect 315818 496170 315888 496226
rect 315568 496102 315888 496170
rect 315568 496046 315638 496102
rect 315694 496046 315762 496102
rect 315818 496046 315888 496102
rect 315568 495978 315888 496046
rect 315568 495922 315638 495978
rect 315694 495922 315762 495978
rect 315818 495922 315888 495978
rect 315568 495888 315888 495922
rect 346288 496350 346608 496384
rect 346288 496294 346358 496350
rect 346414 496294 346482 496350
rect 346538 496294 346608 496350
rect 346288 496226 346608 496294
rect 346288 496170 346358 496226
rect 346414 496170 346482 496226
rect 346538 496170 346608 496226
rect 346288 496102 346608 496170
rect 346288 496046 346358 496102
rect 346414 496046 346482 496102
rect 346538 496046 346608 496102
rect 346288 495978 346608 496046
rect 346288 495922 346358 495978
rect 346414 495922 346482 495978
rect 346538 495922 346608 495978
rect 346288 495888 346608 495922
rect 377008 496350 377328 496384
rect 377008 496294 377078 496350
rect 377134 496294 377202 496350
rect 377258 496294 377328 496350
rect 377008 496226 377328 496294
rect 377008 496170 377078 496226
rect 377134 496170 377202 496226
rect 377258 496170 377328 496226
rect 377008 496102 377328 496170
rect 377008 496046 377078 496102
rect 377134 496046 377202 496102
rect 377258 496046 377328 496102
rect 377008 495978 377328 496046
rect 377008 495922 377078 495978
rect 377134 495922 377202 495978
rect 377258 495922 377328 495978
rect 377008 495888 377328 495922
rect 407728 496350 408048 496384
rect 407728 496294 407798 496350
rect 407854 496294 407922 496350
rect 407978 496294 408048 496350
rect 407728 496226 408048 496294
rect 407728 496170 407798 496226
rect 407854 496170 407922 496226
rect 407978 496170 408048 496226
rect 407728 496102 408048 496170
rect 407728 496046 407798 496102
rect 407854 496046 407922 496102
rect 407978 496046 408048 496102
rect 407728 495978 408048 496046
rect 407728 495922 407798 495978
rect 407854 495922 407922 495978
rect 407978 495922 408048 495978
rect 407728 495888 408048 495922
rect 438448 496350 438768 496384
rect 438448 496294 438518 496350
rect 438574 496294 438642 496350
rect 438698 496294 438768 496350
rect 438448 496226 438768 496294
rect 438448 496170 438518 496226
rect 438574 496170 438642 496226
rect 438698 496170 438768 496226
rect 438448 496102 438768 496170
rect 438448 496046 438518 496102
rect 438574 496046 438642 496102
rect 438698 496046 438768 496102
rect 438448 495978 438768 496046
rect 438448 495922 438518 495978
rect 438574 495922 438642 495978
rect 438698 495922 438768 495978
rect 438448 495888 438768 495922
rect 469168 496350 469488 496384
rect 469168 496294 469238 496350
rect 469294 496294 469362 496350
rect 469418 496294 469488 496350
rect 469168 496226 469488 496294
rect 469168 496170 469238 496226
rect 469294 496170 469362 496226
rect 469418 496170 469488 496226
rect 469168 496102 469488 496170
rect 469168 496046 469238 496102
rect 469294 496046 469362 496102
rect 469418 496046 469488 496102
rect 469168 495978 469488 496046
rect 469168 495922 469238 495978
rect 469294 495922 469362 495978
rect 469418 495922 469488 495978
rect 469168 495888 469488 495922
rect 499888 496350 500208 496384
rect 499888 496294 499958 496350
rect 500014 496294 500082 496350
rect 500138 496294 500208 496350
rect 499888 496226 500208 496294
rect 499888 496170 499958 496226
rect 500014 496170 500082 496226
rect 500138 496170 500208 496226
rect 499888 496102 500208 496170
rect 499888 496046 499958 496102
rect 500014 496046 500082 496102
rect 500138 496046 500208 496102
rect 499888 495978 500208 496046
rect 499888 495922 499958 495978
rect 500014 495922 500082 495978
rect 500138 495922 500208 495978
rect 499888 495888 500208 495922
rect 530608 496350 530928 496384
rect 530608 496294 530678 496350
rect 530734 496294 530802 496350
rect 530858 496294 530928 496350
rect 530608 496226 530928 496294
rect 530608 496170 530678 496226
rect 530734 496170 530802 496226
rect 530858 496170 530928 496226
rect 530608 496102 530928 496170
rect 530608 496046 530678 496102
rect 530734 496046 530802 496102
rect 530858 496046 530928 496102
rect 530608 495978 530928 496046
rect 530608 495922 530678 495978
rect 530734 495922 530802 495978
rect 530858 495922 530928 495978
rect 530608 495888 530928 495922
rect 111154 490294 111250 490350
rect 111306 490294 111374 490350
rect 111430 490294 111498 490350
rect 111554 490294 111622 490350
rect 111678 490294 111774 490350
rect 111154 490226 111774 490294
rect 111154 490170 111250 490226
rect 111306 490170 111374 490226
rect 111430 490170 111498 490226
rect 111554 490170 111622 490226
rect 111678 490170 111774 490226
rect 111154 490102 111774 490170
rect 111154 490046 111250 490102
rect 111306 490046 111374 490102
rect 111430 490046 111498 490102
rect 111554 490046 111622 490102
rect 111678 490046 111774 490102
rect 111154 489978 111774 490046
rect 111154 489922 111250 489978
rect 111306 489922 111374 489978
rect 111430 489922 111498 489978
rect 111554 489922 111622 489978
rect 111678 489922 111774 489978
rect 96874 478294 96970 478350
rect 97026 478294 97094 478350
rect 97150 478294 97218 478350
rect 97274 478294 97342 478350
rect 97398 478294 97494 478350
rect 96874 478226 97494 478294
rect 96874 478170 96970 478226
rect 97026 478170 97094 478226
rect 97150 478170 97218 478226
rect 97274 478170 97342 478226
rect 97398 478170 97494 478226
rect 96874 478102 97494 478170
rect 96874 478046 96970 478102
rect 97026 478046 97094 478102
rect 97150 478046 97218 478102
rect 97274 478046 97342 478102
rect 97398 478046 97494 478102
rect 96874 477978 97494 478046
rect 96874 477922 96970 477978
rect 97026 477922 97094 477978
rect 97150 477922 97218 477978
rect 97274 477922 97342 477978
rect 97398 477922 97494 477978
rect 96874 460350 97494 477922
rect 100528 478350 100848 478384
rect 100528 478294 100598 478350
rect 100654 478294 100722 478350
rect 100778 478294 100848 478350
rect 100528 478226 100848 478294
rect 100528 478170 100598 478226
rect 100654 478170 100722 478226
rect 100778 478170 100848 478226
rect 100528 478102 100848 478170
rect 100528 478046 100598 478102
rect 100654 478046 100722 478102
rect 100778 478046 100848 478102
rect 100528 477978 100848 478046
rect 100528 477922 100598 477978
rect 100654 477922 100722 477978
rect 100778 477922 100848 477978
rect 100528 477888 100848 477922
rect 111154 472350 111774 489922
rect 115888 490350 116208 490384
rect 115888 490294 115958 490350
rect 116014 490294 116082 490350
rect 116138 490294 116208 490350
rect 115888 490226 116208 490294
rect 115888 490170 115958 490226
rect 116014 490170 116082 490226
rect 116138 490170 116208 490226
rect 115888 490102 116208 490170
rect 115888 490046 115958 490102
rect 116014 490046 116082 490102
rect 116138 490046 116208 490102
rect 115888 489978 116208 490046
rect 115888 489922 115958 489978
rect 116014 489922 116082 489978
rect 116138 489922 116208 489978
rect 115888 489888 116208 489922
rect 146608 490350 146928 490384
rect 146608 490294 146678 490350
rect 146734 490294 146802 490350
rect 146858 490294 146928 490350
rect 146608 490226 146928 490294
rect 146608 490170 146678 490226
rect 146734 490170 146802 490226
rect 146858 490170 146928 490226
rect 146608 490102 146928 490170
rect 146608 490046 146678 490102
rect 146734 490046 146802 490102
rect 146858 490046 146928 490102
rect 146608 489978 146928 490046
rect 146608 489922 146678 489978
rect 146734 489922 146802 489978
rect 146858 489922 146928 489978
rect 146608 489888 146928 489922
rect 177328 490350 177648 490384
rect 177328 490294 177398 490350
rect 177454 490294 177522 490350
rect 177578 490294 177648 490350
rect 177328 490226 177648 490294
rect 177328 490170 177398 490226
rect 177454 490170 177522 490226
rect 177578 490170 177648 490226
rect 177328 490102 177648 490170
rect 177328 490046 177398 490102
rect 177454 490046 177522 490102
rect 177578 490046 177648 490102
rect 177328 489978 177648 490046
rect 177328 489922 177398 489978
rect 177454 489922 177522 489978
rect 177578 489922 177648 489978
rect 177328 489888 177648 489922
rect 208048 490350 208368 490384
rect 208048 490294 208118 490350
rect 208174 490294 208242 490350
rect 208298 490294 208368 490350
rect 208048 490226 208368 490294
rect 208048 490170 208118 490226
rect 208174 490170 208242 490226
rect 208298 490170 208368 490226
rect 208048 490102 208368 490170
rect 208048 490046 208118 490102
rect 208174 490046 208242 490102
rect 208298 490046 208368 490102
rect 208048 489978 208368 490046
rect 208048 489922 208118 489978
rect 208174 489922 208242 489978
rect 208298 489922 208368 489978
rect 208048 489888 208368 489922
rect 238768 490350 239088 490384
rect 238768 490294 238838 490350
rect 238894 490294 238962 490350
rect 239018 490294 239088 490350
rect 238768 490226 239088 490294
rect 238768 490170 238838 490226
rect 238894 490170 238962 490226
rect 239018 490170 239088 490226
rect 238768 490102 239088 490170
rect 238768 490046 238838 490102
rect 238894 490046 238962 490102
rect 239018 490046 239088 490102
rect 238768 489978 239088 490046
rect 238768 489922 238838 489978
rect 238894 489922 238962 489978
rect 239018 489922 239088 489978
rect 238768 489888 239088 489922
rect 269488 490350 269808 490384
rect 269488 490294 269558 490350
rect 269614 490294 269682 490350
rect 269738 490294 269808 490350
rect 269488 490226 269808 490294
rect 269488 490170 269558 490226
rect 269614 490170 269682 490226
rect 269738 490170 269808 490226
rect 269488 490102 269808 490170
rect 269488 490046 269558 490102
rect 269614 490046 269682 490102
rect 269738 490046 269808 490102
rect 269488 489978 269808 490046
rect 269488 489922 269558 489978
rect 269614 489922 269682 489978
rect 269738 489922 269808 489978
rect 269488 489888 269808 489922
rect 300208 490350 300528 490384
rect 300208 490294 300278 490350
rect 300334 490294 300402 490350
rect 300458 490294 300528 490350
rect 300208 490226 300528 490294
rect 300208 490170 300278 490226
rect 300334 490170 300402 490226
rect 300458 490170 300528 490226
rect 300208 490102 300528 490170
rect 300208 490046 300278 490102
rect 300334 490046 300402 490102
rect 300458 490046 300528 490102
rect 300208 489978 300528 490046
rect 300208 489922 300278 489978
rect 300334 489922 300402 489978
rect 300458 489922 300528 489978
rect 300208 489888 300528 489922
rect 330928 490350 331248 490384
rect 330928 490294 330998 490350
rect 331054 490294 331122 490350
rect 331178 490294 331248 490350
rect 330928 490226 331248 490294
rect 330928 490170 330998 490226
rect 331054 490170 331122 490226
rect 331178 490170 331248 490226
rect 330928 490102 331248 490170
rect 330928 490046 330998 490102
rect 331054 490046 331122 490102
rect 331178 490046 331248 490102
rect 330928 489978 331248 490046
rect 330928 489922 330998 489978
rect 331054 489922 331122 489978
rect 331178 489922 331248 489978
rect 330928 489888 331248 489922
rect 361648 490350 361968 490384
rect 361648 490294 361718 490350
rect 361774 490294 361842 490350
rect 361898 490294 361968 490350
rect 361648 490226 361968 490294
rect 361648 490170 361718 490226
rect 361774 490170 361842 490226
rect 361898 490170 361968 490226
rect 361648 490102 361968 490170
rect 361648 490046 361718 490102
rect 361774 490046 361842 490102
rect 361898 490046 361968 490102
rect 361648 489978 361968 490046
rect 361648 489922 361718 489978
rect 361774 489922 361842 489978
rect 361898 489922 361968 489978
rect 361648 489888 361968 489922
rect 392368 490350 392688 490384
rect 392368 490294 392438 490350
rect 392494 490294 392562 490350
rect 392618 490294 392688 490350
rect 392368 490226 392688 490294
rect 392368 490170 392438 490226
rect 392494 490170 392562 490226
rect 392618 490170 392688 490226
rect 392368 490102 392688 490170
rect 392368 490046 392438 490102
rect 392494 490046 392562 490102
rect 392618 490046 392688 490102
rect 392368 489978 392688 490046
rect 392368 489922 392438 489978
rect 392494 489922 392562 489978
rect 392618 489922 392688 489978
rect 392368 489888 392688 489922
rect 423088 490350 423408 490384
rect 423088 490294 423158 490350
rect 423214 490294 423282 490350
rect 423338 490294 423408 490350
rect 423088 490226 423408 490294
rect 423088 490170 423158 490226
rect 423214 490170 423282 490226
rect 423338 490170 423408 490226
rect 423088 490102 423408 490170
rect 423088 490046 423158 490102
rect 423214 490046 423282 490102
rect 423338 490046 423408 490102
rect 423088 489978 423408 490046
rect 423088 489922 423158 489978
rect 423214 489922 423282 489978
rect 423338 489922 423408 489978
rect 423088 489888 423408 489922
rect 453808 490350 454128 490384
rect 453808 490294 453878 490350
rect 453934 490294 454002 490350
rect 454058 490294 454128 490350
rect 453808 490226 454128 490294
rect 453808 490170 453878 490226
rect 453934 490170 454002 490226
rect 454058 490170 454128 490226
rect 453808 490102 454128 490170
rect 453808 490046 453878 490102
rect 453934 490046 454002 490102
rect 454058 490046 454128 490102
rect 453808 489978 454128 490046
rect 453808 489922 453878 489978
rect 453934 489922 454002 489978
rect 454058 489922 454128 489978
rect 453808 489888 454128 489922
rect 484528 490350 484848 490384
rect 484528 490294 484598 490350
rect 484654 490294 484722 490350
rect 484778 490294 484848 490350
rect 484528 490226 484848 490294
rect 484528 490170 484598 490226
rect 484654 490170 484722 490226
rect 484778 490170 484848 490226
rect 484528 490102 484848 490170
rect 484528 490046 484598 490102
rect 484654 490046 484722 490102
rect 484778 490046 484848 490102
rect 484528 489978 484848 490046
rect 484528 489922 484598 489978
rect 484654 489922 484722 489978
rect 484778 489922 484848 489978
rect 484528 489888 484848 489922
rect 515248 490350 515568 490384
rect 515248 490294 515318 490350
rect 515374 490294 515442 490350
rect 515498 490294 515568 490350
rect 515248 490226 515568 490294
rect 515248 490170 515318 490226
rect 515374 490170 515442 490226
rect 515498 490170 515568 490226
rect 515248 490102 515568 490170
rect 515248 490046 515318 490102
rect 515374 490046 515442 490102
rect 515498 490046 515568 490102
rect 515248 489978 515568 490046
rect 515248 489922 515318 489978
rect 515374 489922 515442 489978
rect 515498 489922 515568 489978
rect 515248 489888 515568 489922
rect 545968 490350 546288 490384
rect 545968 490294 546038 490350
rect 546094 490294 546162 490350
rect 546218 490294 546288 490350
rect 545968 490226 546288 490294
rect 545968 490170 546038 490226
rect 546094 490170 546162 490226
rect 546218 490170 546288 490226
rect 545968 490102 546288 490170
rect 545968 490046 546038 490102
rect 546094 490046 546162 490102
rect 546218 490046 546288 490102
rect 545968 489978 546288 490046
rect 545968 489922 546038 489978
rect 546094 489922 546162 489978
rect 546218 489922 546288 489978
rect 545968 489888 546288 489922
rect 561154 490350 561774 507922
rect 561154 490294 561250 490350
rect 561306 490294 561374 490350
rect 561430 490294 561498 490350
rect 561554 490294 561622 490350
rect 561678 490294 561774 490350
rect 561154 490226 561774 490294
rect 561154 490170 561250 490226
rect 561306 490170 561374 490226
rect 561430 490170 561498 490226
rect 561554 490170 561622 490226
rect 561678 490170 561774 490226
rect 561154 490102 561774 490170
rect 561154 490046 561250 490102
rect 561306 490046 561374 490102
rect 561430 490046 561498 490102
rect 561554 490046 561622 490102
rect 561678 490046 561774 490102
rect 561154 489978 561774 490046
rect 561154 489922 561250 489978
rect 561306 489922 561374 489978
rect 561430 489922 561498 489978
rect 561554 489922 561622 489978
rect 561678 489922 561774 489978
rect 131248 478350 131568 478384
rect 131248 478294 131318 478350
rect 131374 478294 131442 478350
rect 131498 478294 131568 478350
rect 131248 478226 131568 478294
rect 131248 478170 131318 478226
rect 131374 478170 131442 478226
rect 131498 478170 131568 478226
rect 131248 478102 131568 478170
rect 131248 478046 131318 478102
rect 131374 478046 131442 478102
rect 131498 478046 131568 478102
rect 131248 477978 131568 478046
rect 131248 477922 131318 477978
rect 131374 477922 131442 477978
rect 131498 477922 131568 477978
rect 131248 477888 131568 477922
rect 161968 478350 162288 478384
rect 161968 478294 162038 478350
rect 162094 478294 162162 478350
rect 162218 478294 162288 478350
rect 161968 478226 162288 478294
rect 161968 478170 162038 478226
rect 162094 478170 162162 478226
rect 162218 478170 162288 478226
rect 161968 478102 162288 478170
rect 161968 478046 162038 478102
rect 162094 478046 162162 478102
rect 162218 478046 162288 478102
rect 161968 477978 162288 478046
rect 161968 477922 162038 477978
rect 162094 477922 162162 477978
rect 162218 477922 162288 477978
rect 161968 477888 162288 477922
rect 192688 478350 193008 478384
rect 192688 478294 192758 478350
rect 192814 478294 192882 478350
rect 192938 478294 193008 478350
rect 192688 478226 193008 478294
rect 192688 478170 192758 478226
rect 192814 478170 192882 478226
rect 192938 478170 193008 478226
rect 192688 478102 193008 478170
rect 192688 478046 192758 478102
rect 192814 478046 192882 478102
rect 192938 478046 193008 478102
rect 192688 477978 193008 478046
rect 192688 477922 192758 477978
rect 192814 477922 192882 477978
rect 192938 477922 193008 477978
rect 192688 477888 193008 477922
rect 223408 478350 223728 478384
rect 223408 478294 223478 478350
rect 223534 478294 223602 478350
rect 223658 478294 223728 478350
rect 223408 478226 223728 478294
rect 223408 478170 223478 478226
rect 223534 478170 223602 478226
rect 223658 478170 223728 478226
rect 223408 478102 223728 478170
rect 223408 478046 223478 478102
rect 223534 478046 223602 478102
rect 223658 478046 223728 478102
rect 223408 477978 223728 478046
rect 223408 477922 223478 477978
rect 223534 477922 223602 477978
rect 223658 477922 223728 477978
rect 223408 477888 223728 477922
rect 254128 478350 254448 478384
rect 254128 478294 254198 478350
rect 254254 478294 254322 478350
rect 254378 478294 254448 478350
rect 254128 478226 254448 478294
rect 254128 478170 254198 478226
rect 254254 478170 254322 478226
rect 254378 478170 254448 478226
rect 254128 478102 254448 478170
rect 254128 478046 254198 478102
rect 254254 478046 254322 478102
rect 254378 478046 254448 478102
rect 254128 477978 254448 478046
rect 254128 477922 254198 477978
rect 254254 477922 254322 477978
rect 254378 477922 254448 477978
rect 254128 477888 254448 477922
rect 284848 478350 285168 478384
rect 284848 478294 284918 478350
rect 284974 478294 285042 478350
rect 285098 478294 285168 478350
rect 284848 478226 285168 478294
rect 284848 478170 284918 478226
rect 284974 478170 285042 478226
rect 285098 478170 285168 478226
rect 284848 478102 285168 478170
rect 284848 478046 284918 478102
rect 284974 478046 285042 478102
rect 285098 478046 285168 478102
rect 284848 477978 285168 478046
rect 284848 477922 284918 477978
rect 284974 477922 285042 477978
rect 285098 477922 285168 477978
rect 284848 477888 285168 477922
rect 315568 478350 315888 478384
rect 315568 478294 315638 478350
rect 315694 478294 315762 478350
rect 315818 478294 315888 478350
rect 315568 478226 315888 478294
rect 315568 478170 315638 478226
rect 315694 478170 315762 478226
rect 315818 478170 315888 478226
rect 315568 478102 315888 478170
rect 315568 478046 315638 478102
rect 315694 478046 315762 478102
rect 315818 478046 315888 478102
rect 315568 477978 315888 478046
rect 315568 477922 315638 477978
rect 315694 477922 315762 477978
rect 315818 477922 315888 477978
rect 315568 477888 315888 477922
rect 346288 478350 346608 478384
rect 346288 478294 346358 478350
rect 346414 478294 346482 478350
rect 346538 478294 346608 478350
rect 346288 478226 346608 478294
rect 346288 478170 346358 478226
rect 346414 478170 346482 478226
rect 346538 478170 346608 478226
rect 346288 478102 346608 478170
rect 346288 478046 346358 478102
rect 346414 478046 346482 478102
rect 346538 478046 346608 478102
rect 346288 477978 346608 478046
rect 346288 477922 346358 477978
rect 346414 477922 346482 477978
rect 346538 477922 346608 477978
rect 346288 477888 346608 477922
rect 377008 478350 377328 478384
rect 377008 478294 377078 478350
rect 377134 478294 377202 478350
rect 377258 478294 377328 478350
rect 377008 478226 377328 478294
rect 377008 478170 377078 478226
rect 377134 478170 377202 478226
rect 377258 478170 377328 478226
rect 377008 478102 377328 478170
rect 377008 478046 377078 478102
rect 377134 478046 377202 478102
rect 377258 478046 377328 478102
rect 377008 477978 377328 478046
rect 377008 477922 377078 477978
rect 377134 477922 377202 477978
rect 377258 477922 377328 477978
rect 377008 477888 377328 477922
rect 407728 478350 408048 478384
rect 407728 478294 407798 478350
rect 407854 478294 407922 478350
rect 407978 478294 408048 478350
rect 407728 478226 408048 478294
rect 407728 478170 407798 478226
rect 407854 478170 407922 478226
rect 407978 478170 408048 478226
rect 407728 478102 408048 478170
rect 407728 478046 407798 478102
rect 407854 478046 407922 478102
rect 407978 478046 408048 478102
rect 407728 477978 408048 478046
rect 407728 477922 407798 477978
rect 407854 477922 407922 477978
rect 407978 477922 408048 477978
rect 407728 477888 408048 477922
rect 438448 478350 438768 478384
rect 438448 478294 438518 478350
rect 438574 478294 438642 478350
rect 438698 478294 438768 478350
rect 438448 478226 438768 478294
rect 438448 478170 438518 478226
rect 438574 478170 438642 478226
rect 438698 478170 438768 478226
rect 438448 478102 438768 478170
rect 438448 478046 438518 478102
rect 438574 478046 438642 478102
rect 438698 478046 438768 478102
rect 438448 477978 438768 478046
rect 438448 477922 438518 477978
rect 438574 477922 438642 477978
rect 438698 477922 438768 477978
rect 438448 477888 438768 477922
rect 469168 478350 469488 478384
rect 469168 478294 469238 478350
rect 469294 478294 469362 478350
rect 469418 478294 469488 478350
rect 469168 478226 469488 478294
rect 469168 478170 469238 478226
rect 469294 478170 469362 478226
rect 469418 478170 469488 478226
rect 469168 478102 469488 478170
rect 469168 478046 469238 478102
rect 469294 478046 469362 478102
rect 469418 478046 469488 478102
rect 469168 477978 469488 478046
rect 469168 477922 469238 477978
rect 469294 477922 469362 477978
rect 469418 477922 469488 477978
rect 469168 477888 469488 477922
rect 499888 478350 500208 478384
rect 499888 478294 499958 478350
rect 500014 478294 500082 478350
rect 500138 478294 500208 478350
rect 499888 478226 500208 478294
rect 499888 478170 499958 478226
rect 500014 478170 500082 478226
rect 500138 478170 500208 478226
rect 499888 478102 500208 478170
rect 499888 478046 499958 478102
rect 500014 478046 500082 478102
rect 500138 478046 500208 478102
rect 499888 477978 500208 478046
rect 499888 477922 499958 477978
rect 500014 477922 500082 477978
rect 500138 477922 500208 477978
rect 499888 477888 500208 477922
rect 530608 478350 530928 478384
rect 530608 478294 530678 478350
rect 530734 478294 530802 478350
rect 530858 478294 530928 478350
rect 530608 478226 530928 478294
rect 530608 478170 530678 478226
rect 530734 478170 530802 478226
rect 530858 478170 530928 478226
rect 530608 478102 530928 478170
rect 530608 478046 530678 478102
rect 530734 478046 530802 478102
rect 530858 478046 530928 478102
rect 530608 477978 530928 478046
rect 530608 477922 530678 477978
rect 530734 477922 530802 477978
rect 530858 477922 530928 477978
rect 530608 477888 530928 477922
rect 111154 472294 111250 472350
rect 111306 472294 111374 472350
rect 111430 472294 111498 472350
rect 111554 472294 111622 472350
rect 111678 472294 111774 472350
rect 111154 472226 111774 472294
rect 111154 472170 111250 472226
rect 111306 472170 111374 472226
rect 111430 472170 111498 472226
rect 111554 472170 111622 472226
rect 111678 472170 111774 472226
rect 111154 472102 111774 472170
rect 111154 472046 111250 472102
rect 111306 472046 111374 472102
rect 111430 472046 111498 472102
rect 111554 472046 111622 472102
rect 111678 472046 111774 472102
rect 111154 471978 111774 472046
rect 111154 471922 111250 471978
rect 111306 471922 111374 471978
rect 111430 471922 111498 471978
rect 111554 471922 111622 471978
rect 111678 471922 111774 471978
rect 96874 460294 96970 460350
rect 97026 460294 97094 460350
rect 97150 460294 97218 460350
rect 97274 460294 97342 460350
rect 97398 460294 97494 460350
rect 96874 460226 97494 460294
rect 96874 460170 96970 460226
rect 97026 460170 97094 460226
rect 97150 460170 97218 460226
rect 97274 460170 97342 460226
rect 97398 460170 97494 460226
rect 96874 460102 97494 460170
rect 96874 460046 96970 460102
rect 97026 460046 97094 460102
rect 97150 460046 97218 460102
rect 97274 460046 97342 460102
rect 97398 460046 97494 460102
rect 96874 459978 97494 460046
rect 96874 459922 96970 459978
rect 97026 459922 97094 459978
rect 97150 459922 97218 459978
rect 97274 459922 97342 459978
rect 97398 459922 97494 459978
rect 96874 442350 97494 459922
rect 100528 460350 100848 460384
rect 100528 460294 100598 460350
rect 100654 460294 100722 460350
rect 100778 460294 100848 460350
rect 100528 460226 100848 460294
rect 100528 460170 100598 460226
rect 100654 460170 100722 460226
rect 100778 460170 100848 460226
rect 100528 460102 100848 460170
rect 100528 460046 100598 460102
rect 100654 460046 100722 460102
rect 100778 460046 100848 460102
rect 100528 459978 100848 460046
rect 100528 459922 100598 459978
rect 100654 459922 100722 459978
rect 100778 459922 100848 459978
rect 100528 459888 100848 459922
rect 111154 454350 111774 471922
rect 115888 472350 116208 472384
rect 115888 472294 115958 472350
rect 116014 472294 116082 472350
rect 116138 472294 116208 472350
rect 115888 472226 116208 472294
rect 115888 472170 115958 472226
rect 116014 472170 116082 472226
rect 116138 472170 116208 472226
rect 115888 472102 116208 472170
rect 115888 472046 115958 472102
rect 116014 472046 116082 472102
rect 116138 472046 116208 472102
rect 115888 471978 116208 472046
rect 115888 471922 115958 471978
rect 116014 471922 116082 471978
rect 116138 471922 116208 471978
rect 115888 471888 116208 471922
rect 146608 472350 146928 472384
rect 146608 472294 146678 472350
rect 146734 472294 146802 472350
rect 146858 472294 146928 472350
rect 146608 472226 146928 472294
rect 146608 472170 146678 472226
rect 146734 472170 146802 472226
rect 146858 472170 146928 472226
rect 146608 472102 146928 472170
rect 146608 472046 146678 472102
rect 146734 472046 146802 472102
rect 146858 472046 146928 472102
rect 146608 471978 146928 472046
rect 146608 471922 146678 471978
rect 146734 471922 146802 471978
rect 146858 471922 146928 471978
rect 146608 471888 146928 471922
rect 177328 472350 177648 472384
rect 177328 472294 177398 472350
rect 177454 472294 177522 472350
rect 177578 472294 177648 472350
rect 177328 472226 177648 472294
rect 177328 472170 177398 472226
rect 177454 472170 177522 472226
rect 177578 472170 177648 472226
rect 177328 472102 177648 472170
rect 177328 472046 177398 472102
rect 177454 472046 177522 472102
rect 177578 472046 177648 472102
rect 177328 471978 177648 472046
rect 177328 471922 177398 471978
rect 177454 471922 177522 471978
rect 177578 471922 177648 471978
rect 177328 471888 177648 471922
rect 208048 472350 208368 472384
rect 208048 472294 208118 472350
rect 208174 472294 208242 472350
rect 208298 472294 208368 472350
rect 208048 472226 208368 472294
rect 208048 472170 208118 472226
rect 208174 472170 208242 472226
rect 208298 472170 208368 472226
rect 208048 472102 208368 472170
rect 208048 472046 208118 472102
rect 208174 472046 208242 472102
rect 208298 472046 208368 472102
rect 208048 471978 208368 472046
rect 208048 471922 208118 471978
rect 208174 471922 208242 471978
rect 208298 471922 208368 471978
rect 208048 471888 208368 471922
rect 238768 472350 239088 472384
rect 238768 472294 238838 472350
rect 238894 472294 238962 472350
rect 239018 472294 239088 472350
rect 238768 472226 239088 472294
rect 238768 472170 238838 472226
rect 238894 472170 238962 472226
rect 239018 472170 239088 472226
rect 238768 472102 239088 472170
rect 238768 472046 238838 472102
rect 238894 472046 238962 472102
rect 239018 472046 239088 472102
rect 238768 471978 239088 472046
rect 238768 471922 238838 471978
rect 238894 471922 238962 471978
rect 239018 471922 239088 471978
rect 238768 471888 239088 471922
rect 269488 472350 269808 472384
rect 269488 472294 269558 472350
rect 269614 472294 269682 472350
rect 269738 472294 269808 472350
rect 269488 472226 269808 472294
rect 269488 472170 269558 472226
rect 269614 472170 269682 472226
rect 269738 472170 269808 472226
rect 269488 472102 269808 472170
rect 269488 472046 269558 472102
rect 269614 472046 269682 472102
rect 269738 472046 269808 472102
rect 269488 471978 269808 472046
rect 269488 471922 269558 471978
rect 269614 471922 269682 471978
rect 269738 471922 269808 471978
rect 269488 471888 269808 471922
rect 300208 472350 300528 472384
rect 300208 472294 300278 472350
rect 300334 472294 300402 472350
rect 300458 472294 300528 472350
rect 300208 472226 300528 472294
rect 300208 472170 300278 472226
rect 300334 472170 300402 472226
rect 300458 472170 300528 472226
rect 300208 472102 300528 472170
rect 300208 472046 300278 472102
rect 300334 472046 300402 472102
rect 300458 472046 300528 472102
rect 300208 471978 300528 472046
rect 300208 471922 300278 471978
rect 300334 471922 300402 471978
rect 300458 471922 300528 471978
rect 300208 471888 300528 471922
rect 330928 472350 331248 472384
rect 330928 472294 330998 472350
rect 331054 472294 331122 472350
rect 331178 472294 331248 472350
rect 330928 472226 331248 472294
rect 330928 472170 330998 472226
rect 331054 472170 331122 472226
rect 331178 472170 331248 472226
rect 330928 472102 331248 472170
rect 330928 472046 330998 472102
rect 331054 472046 331122 472102
rect 331178 472046 331248 472102
rect 330928 471978 331248 472046
rect 330928 471922 330998 471978
rect 331054 471922 331122 471978
rect 331178 471922 331248 471978
rect 330928 471888 331248 471922
rect 361648 472350 361968 472384
rect 361648 472294 361718 472350
rect 361774 472294 361842 472350
rect 361898 472294 361968 472350
rect 361648 472226 361968 472294
rect 361648 472170 361718 472226
rect 361774 472170 361842 472226
rect 361898 472170 361968 472226
rect 361648 472102 361968 472170
rect 361648 472046 361718 472102
rect 361774 472046 361842 472102
rect 361898 472046 361968 472102
rect 361648 471978 361968 472046
rect 361648 471922 361718 471978
rect 361774 471922 361842 471978
rect 361898 471922 361968 471978
rect 361648 471888 361968 471922
rect 392368 472350 392688 472384
rect 392368 472294 392438 472350
rect 392494 472294 392562 472350
rect 392618 472294 392688 472350
rect 392368 472226 392688 472294
rect 392368 472170 392438 472226
rect 392494 472170 392562 472226
rect 392618 472170 392688 472226
rect 392368 472102 392688 472170
rect 392368 472046 392438 472102
rect 392494 472046 392562 472102
rect 392618 472046 392688 472102
rect 392368 471978 392688 472046
rect 392368 471922 392438 471978
rect 392494 471922 392562 471978
rect 392618 471922 392688 471978
rect 392368 471888 392688 471922
rect 423088 472350 423408 472384
rect 423088 472294 423158 472350
rect 423214 472294 423282 472350
rect 423338 472294 423408 472350
rect 423088 472226 423408 472294
rect 423088 472170 423158 472226
rect 423214 472170 423282 472226
rect 423338 472170 423408 472226
rect 423088 472102 423408 472170
rect 423088 472046 423158 472102
rect 423214 472046 423282 472102
rect 423338 472046 423408 472102
rect 423088 471978 423408 472046
rect 423088 471922 423158 471978
rect 423214 471922 423282 471978
rect 423338 471922 423408 471978
rect 423088 471888 423408 471922
rect 453808 472350 454128 472384
rect 453808 472294 453878 472350
rect 453934 472294 454002 472350
rect 454058 472294 454128 472350
rect 453808 472226 454128 472294
rect 453808 472170 453878 472226
rect 453934 472170 454002 472226
rect 454058 472170 454128 472226
rect 453808 472102 454128 472170
rect 453808 472046 453878 472102
rect 453934 472046 454002 472102
rect 454058 472046 454128 472102
rect 453808 471978 454128 472046
rect 453808 471922 453878 471978
rect 453934 471922 454002 471978
rect 454058 471922 454128 471978
rect 453808 471888 454128 471922
rect 484528 472350 484848 472384
rect 484528 472294 484598 472350
rect 484654 472294 484722 472350
rect 484778 472294 484848 472350
rect 484528 472226 484848 472294
rect 484528 472170 484598 472226
rect 484654 472170 484722 472226
rect 484778 472170 484848 472226
rect 484528 472102 484848 472170
rect 484528 472046 484598 472102
rect 484654 472046 484722 472102
rect 484778 472046 484848 472102
rect 484528 471978 484848 472046
rect 484528 471922 484598 471978
rect 484654 471922 484722 471978
rect 484778 471922 484848 471978
rect 484528 471888 484848 471922
rect 515248 472350 515568 472384
rect 515248 472294 515318 472350
rect 515374 472294 515442 472350
rect 515498 472294 515568 472350
rect 515248 472226 515568 472294
rect 515248 472170 515318 472226
rect 515374 472170 515442 472226
rect 515498 472170 515568 472226
rect 515248 472102 515568 472170
rect 515248 472046 515318 472102
rect 515374 472046 515442 472102
rect 515498 472046 515568 472102
rect 515248 471978 515568 472046
rect 515248 471922 515318 471978
rect 515374 471922 515442 471978
rect 515498 471922 515568 471978
rect 515248 471888 515568 471922
rect 545968 472350 546288 472384
rect 545968 472294 546038 472350
rect 546094 472294 546162 472350
rect 546218 472294 546288 472350
rect 545968 472226 546288 472294
rect 545968 472170 546038 472226
rect 546094 472170 546162 472226
rect 546218 472170 546288 472226
rect 545968 472102 546288 472170
rect 545968 472046 546038 472102
rect 546094 472046 546162 472102
rect 546218 472046 546288 472102
rect 545968 471978 546288 472046
rect 545968 471922 546038 471978
rect 546094 471922 546162 471978
rect 546218 471922 546288 471978
rect 545968 471888 546288 471922
rect 561154 472350 561774 489922
rect 561154 472294 561250 472350
rect 561306 472294 561374 472350
rect 561430 472294 561498 472350
rect 561554 472294 561622 472350
rect 561678 472294 561774 472350
rect 561154 472226 561774 472294
rect 561154 472170 561250 472226
rect 561306 472170 561374 472226
rect 561430 472170 561498 472226
rect 561554 472170 561622 472226
rect 561678 472170 561774 472226
rect 561154 472102 561774 472170
rect 561154 472046 561250 472102
rect 561306 472046 561374 472102
rect 561430 472046 561498 472102
rect 561554 472046 561622 472102
rect 561678 472046 561774 472102
rect 561154 471978 561774 472046
rect 561154 471922 561250 471978
rect 561306 471922 561374 471978
rect 561430 471922 561498 471978
rect 561554 471922 561622 471978
rect 561678 471922 561774 471978
rect 131248 460350 131568 460384
rect 131248 460294 131318 460350
rect 131374 460294 131442 460350
rect 131498 460294 131568 460350
rect 131248 460226 131568 460294
rect 131248 460170 131318 460226
rect 131374 460170 131442 460226
rect 131498 460170 131568 460226
rect 131248 460102 131568 460170
rect 131248 460046 131318 460102
rect 131374 460046 131442 460102
rect 131498 460046 131568 460102
rect 131248 459978 131568 460046
rect 131248 459922 131318 459978
rect 131374 459922 131442 459978
rect 131498 459922 131568 459978
rect 131248 459888 131568 459922
rect 161968 460350 162288 460384
rect 161968 460294 162038 460350
rect 162094 460294 162162 460350
rect 162218 460294 162288 460350
rect 161968 460226 162288 460294
rect 161968 460170 162038 460226
rect 162094 460170 162162 460226
rect 162218 460170 162288 460226
rect 161968 460102 162288 460170
rect 161968 460046 162038 460102
rect 162094 460046 162162 460102
rect 162218 460046 162288 460102
rect 161968 459978 162288 460046
rect 161968 459922 162038 459978
rect 162094 459922 162162 459978
rect 162218 459922 162288 459978
rect 161968 459888 162288 459922
rect 192688 460350 193008 460384
rect 192688 460294 192758 460350
rect 192814 460294 192882 460350
rect 192938 460294 193008 460350
rect 192688 460226 193008 460294
rect 192688 460170 192758 460226
rect 192814 460170 192882 460226
rect 192938 460170 193008 460226
rect 192688 460102 193008 460170
rect 192688 460046 192758 460102
rect 192814 460046 192882 460102
rect 192938 460046 193008 460102
rect 192688 459978 193008 460046
rect 192688 459922 192758 459978
rect 192814 459922 192882 459978
rect 192938 459922 193008 459978
rect 192688 459888 193008 459922
rect 223408 460350 223728 460384
rect 223408 460294 223478 460350
rect 223534 460294 223602 460350
rect 223658 460294 223728 460350
rect 223408 460226 223728 460294
rect 223408 460170 223478 460226
rect 223534 460170 223602 460226
rect 223658 460170 223728 460226
rect 223408 460102 223728 460170
rect 223408 460046 223478 460102
rect 223534 460046 223602 460102
rect 223658 460046 223728 460102
rect 223408 459978 223728 460046
rect 223408 459922 223478 459978
rect 223534 459922 223602 459978
rect 223658 459922 223728 459978
rect 223408 459888 223728 459922
rect 254128 460350 254448 460384
rect 254128 460294 254198 460350
rect 254254 460294 254322 460350
rect 254378 460294 254448 460350
rect 254128 460226 254448 460294
rect 254128 460170 254198 460226
rect 254254 460170 254322 460226
rect 254378 460170 254448 460226
rect 254128 460102 254448 460170
rect 254128 460046 254198 460102
rect 254254 460046 254322 460102
rect 254378 460046 254448 460102
rect 254128 459978 254448 460046
rect 254128 459922 254198 459978
rect 254254 459922 254322 459978
rect 254378 459922 254448 459978
rect 254128 459888 254448 459922
rect 284848 460350 285168 460384
rect 284848 460294 284918 460350
rect 284974 460294 285042 460350
rect 285098 460294 285168 460350
rect 284848 460226 285168 460294
rect 284848 460170 284918 460226
rect 284974 460170 285042 460226
rect 285098 460170 285168 460226
rect 284848 460102 285168 460170
rect 284848 460046 284918 460102
rect 284974 460046 285042 460102
rect 285098 460046 285168 460102
rect 284848 459978 285168 460046
rect 284848 459922 284918 459978
rect 284974 459922 285042 459978
rect 285098 459922 285168 459978
rect 284848 459888 285168 459922
rect 315568 460350 315888 460384
rect 315568 460294 315638 460350
rect 315694 460294 315762 460350
rect 315818 460294 315888 460350
rect 315568 460226 315888 460294
rect 315568 460170 315638 460226
rect 315694 460170 315762 460226
rect 315818 460170 315888 460226
rect 315568 460102 315888 460170
rect 315568 460046 315638 460102
rect 315694 460046 315762 460102
rect 315818 460046 315888 460102
rect 315568 459978 315888 460046
rect 315568 459922 315638 459978
rect 315694 459922 315762 459978
rect 315818 459922 315888 459978
rect 315568 459888 315888 459922
rect 346288 460350 346608 460384
rect 346288 460294 346358 460350
rect 346414 460294 346482 460350
rect 346538 460294 346608 460350
rect 346288 460226 346608 460294
rect 346288 460170 346358 460226
rect 346414 460170 346482 460226
rect 346538 460170 346608 460226
rect 346288 460102 346608 460170
rect 346288 460046 346358 460102
rect 346414 460046 346482 460102
rect 346538 460046 346608 460102
rect 346288 459978 346608 460046
rect 346288 459922 346358 459978
rect 346414 459922 346482 459978
rect 346538 459922 346608 459978
rect 346288 459888 346608 459922
rect 377008 460350 377328 460384
rect 377008 460294 377078 460350
rect 377134 460294 377202 460350
rect 377258 460294 377328 460350
rect 377008 460226 377328 460294
rect 377008 460170 377078 460226
rect 377134 460170 377202 460226
rect 377258 460170 377328 460226
rect 377008 460102 377328 460170
rect 377008 460046 377078 460102
rect 377134 460046 377202 460102
rect 377258 460046 377328 460102
rect 377008 459978 377328 460046
rect 377008 459922 377078 459978
rect 377134 459922 377202 459978
rect 377258 459922 377328 459978
rect 377008 459888 377328 459922
rect 407728 460350 408048 460384
rect 407728 460294 407798 460350
rect 407854 460294 407922 460350
rect 407978 460294 408048 460350
rect 407728 460226 408048 460294
rect 407728 460170 407798 460226
rect 407854 460170 407922 460226
rect 407978 460170 408048 460226
rect 407728 460102 408048 460170
rect 407728 460046 407798 460102
rect 407854 460046 407922 460102
rect 407978 460046 408048 460102
rect 407728 459978 408048 460046
rect 407728 459922 407798 459978
rect 407854 459922 407922 459978
rect 407978 459922 408048 459978
rect 407728 459888 408048 459922
rect 438448 460350 438768 460384
rect 438448 460294 438518 460350
rect 438574 460294 438642 460350
rect 438698 460294 438768 460350
rect 438448 460226 438768 460294
rect 438448 460170 438518 460226
rect 438574 460170 438642 460226
rect 438698 460170 438768 460226
rect 438448 460102 438768 460170
rect 438448 460046 438518 460102
rect 438574 460046 438642 460102
rect 438698 460046 438768 460102
rect 438448 459978 438768 460046
rect 438448 459922 438518 459978
rect 438574 459922 438642 459978
rect 438698 459922 438768 459978
rect 438448 459888 438768 459922
rect 469168 460350 469488 460384
rect 469168 460294 469238 460350
rect 469294 460294 469362 460350
rect 469418 460294 469488 460350
rect 469168 460226 469488 460294
rect 469168 460170 469238 460226
rect 469294 460170 469362 460226
rect 469418 460170 469488 460226
rect 469168 460102 469488 460170
rect 469168 460046 469238 460102
rect 469294 460046 469362 460102
rect 469418 460046 469488 460102
rect 469168 459978 469488 460046
rect 469168 459922 469238 459978
rect 469294 459922 469362 459978
rect 469418 459922 469488 459978
rect 469168 459888 469488 459922
rect 499888 460350 500208 460384
rect 499888 460294 499958 460350
rect 500014 460294 500082 460350
rect 500138 460294 500208 460350
rect 499888 460226 500208 460294
rect 499888 460170 499958 460226
rect 500014 460170 500082 460226
rect 500138 460170 500208 460226
rect 499888 460102 500208 460170
rect 499888 460046 499958 460102
rect 500014 460046 500082 460102
rect 500138 460046 500208 460102
rect 499888 459978 500208 460046
rect 499888 459922 499958 459978
rect 500014 459922 500082 459978
rect 500138 459922 500208 459978
rect 499888 459888 500208 459922
rect 530608 460350 530928 460384
rect 530608 460294 530678 460350
rect 530734 460294 530802 460350
rect 530858 460294 530928 460350
rect 530608 460226 530928 460294
rect 530608 460170 530678 460226
rect 530734 460170 530802 460226
rect 530858 460170 530928 460226
rect 530608 460102 530928 460170
rect 530608 460046 530678 460102
rect 530734 460046 530802 460102
rect 530858 460046 530928 460102
rect 530608 459978 530928 460046
rect 530608 459922 530678 459978
rect 530734 459922 530802 459978
rect 530858 459922 530928 459978
rect 530608 459888 530928 459922
rect 111154 454294 111250 454350
rect 111306 454294 111374 454350
rect 111430 454294 111498 454350
rect 111554 454294 111622 454350
rect 111678 454294 111774 454350
rect 111154 454226 111774 454294
rect 111154 454170 111250 454226
rect 111306 454170 111374 454226
rect 111430 454170 111498 454226
rect 111554 454170 111622 454226
rect 111678 454170 111774 454226
rect 111154 454102 111774 454170
rect 111154 454046 111250 454102
rect 111306 454046 111374 454102
rect 111430 454046 111498 454102
rect 111554 454046 111622 454102
rect 111678 454046 111774 454102
rect 111154 453978 111774 454046
rect 111154 453922 111250 453978
rect 111306 453922 111374 453978
rect 111430 453922 111498 453978
rect 111554 453922 111622 453978
rect 111678 453922 111774 453978
rect 96874 442294 96970 442350
rect 97026 442294 97094 442350
rect 97150 442294 97218 442350
rect 97274 442294 97342 442350
rect 97398 442294 97494 442350
rect 96874 442226 97494 442294
rect 96874 442170 96970 442226
rect 97026 442170 97094 442226
rect 97150 442170 97218 442226
rect 97274 442170 97342 442226
rect 97398 442170 97494 442226
rect 96874 442102 97494 442170
rect 96874 442046 96970 442102
rect 97026 442046 97094 442102
rect 97150 442046 97218 442102
rect 97274 442046 97342 442102
rect 97398 442046 97494 442102
rect 96874 441978 97494 442046
rect 96874 441922 96970 441978
rect 97026 441922 97094 441978
rect 97150 441922 97218 441978
rect 97274 441922 97342 441978
rect 97398 441922 97494 441978
rect 96874 424350 97494 441922
rect 100528 442350 100848 442384
rect 100528 442294 100598 442350
rect 100654 442294 100722 442350
rect 100778 442294 100848 442350
rect 100528 442226 100848 442294
rect 100528 442170 100598 442226
rect 100654 442170 100722 442226
rect 100778 442170 100848 442226
rect 100528 442102 100848 442170
rect 100528 442046 100598 442102
rect 100654 442046 100722 442102
rect 100778 442046 100848 442102
rect 100528 441978 100848 442046
rect 100528 441922 100598 441978
rect 100654 441922 100722 441978
rect 100778 441922 100848 441978
rect 100528 441888 100848 441922
rect 111154 436350 111774 453922
rect 115888 454350 116208 454384
rect 115888 454294 115958 454350
rect 116014 454294 116082 454350
rect 116138 454294 116208 454350
rect 115888 454226 116208 454294
rect 115888 454170 115958 454226
rect 116014 454170 116082 454226
rect 116138 454170 116208 454226
rect 115888 454102 116208 454170
rect 115888 454046 115958 454102
rect 116014 454046 116082 454102
rect 116138 454046 116208 454102
rect 115888 453978 116208 454046
rect 115888 453922 115958 453978
rect 116014 453922 116082 453978
rect 116138 453922 116208 453978
rect 115888 453888 116208 453922
rect 146608 454350 146928 454384
rect 146608 454294 146678 454350
rect 146734 454294 146802 454350
rect 146858 454294 146928 454350
rect 146608 454226 146928 454294
rect 146608 454170 146678 454226
rect 146734 454170 146802 454226
rect 146858 454170 146928 454226
rect 146608 454102 146928 454170
rect 146608 454046 146678 454102
rect 146734 454046 146802 454102
rect 146858 454046 146928 454102
rect 146608 453978 146928 454046
rect 146608 453922 146678 453978
rect 146734 453922 146802 453978
rect 146858 453922 146928 453978
rect 146608 453888 146928 453922
rect 177328 454350 177648 454384
rect 177328 454294 177398 454350
rect 177454 454294 177522 454350
rect 177578 454294 177648 454350
rect 177328 454226 177648 454294
rect 177328 454170 177398 454226
rect 177454 454170 177522 454226
rect 177578 454170 177648 454226
rect 177328 454102 177648 454170
rect 177328 454046 177398 454102
rect 177454 454046 177522 454102
rect 177578 454046 177648 454102
rect 177328 453978 177648 454046
rect 177328 453922 177398 453978
rect 177454 453922 177522 453978
rect 177578 453922 177648 453978
rect 177328 453888 177648 453922
rect 208048 454350 208368 454384
rect 208048 454294 208118 454350
rect 208174 454294 208242 454350
rect 208298 454294 208368 454350
rect 208048 454226 208368 454294
rect 208048 454170 208118 454226
rect 208174 454170 208242 454226
rect 208298 454170 208368 454226
rect 208048 454102 208368 454170
rect 208048 454046 208118 454102
rect 208174 454046 208242 454102
rect 208298 454046 208368 454102
rect 208048 453978 208368 454046
rect 208048 453922 208118 453978
rect 208174 453922 208242 453978
rect 208298 453922 208368 453978
rect 208048 453888 208368 453922
rect 238768 454350 239088 454384
rect 238768 454294 238838 454350
rect 238894 454294 238962 454350
rect 239018 454294 239088 454350
rect 238768 454226 239088 454294
rect 238768 454170 238838 454226
rect 238894 454170 238962 454226
rect 239018 454170 239088 454226
rect 238768 454102 239088 454170
rect 238768 454046 238838 454102
rect 238894 454046 238962 454102
rect 239018 454046 239088 454102
rect 238768 453978 239088 454046
rect 238768 453922 238838 453978
rect 238894 453922 238962 453978
rect 239018 453922 239088 453978
rect 238768 453888 239088 453922
rect 269488 454350 269808 454384
rect 269488 454294 269558 454350
rect 269614 454294 269682 454350
rect 269738 454294 269808 454350
rect 269488 454226 269808 454294
rect 269488 454170 269558 454226
rect 269614 454170 269682 454226
rect 269738 454170 269808 454226
rect 269488 454102 269808 454170
rect 269488 454046 269558 454102
rect 269614 454046 269682 454102
rect 269738 454046 269808 454102
rect 269488 453978 269808 454046
rect 269488 453922 269558 453978
rect 269614 453922 269682 453978
rect 269738 453922 269808 453978
rect 269488 453888 269808 453922
rect 300208 454350 300528 454384
rect 300208 454294 300278 454350
rect 300334 454294 300402 454350
rect 300458 454294 300528 454350
rect 300208 454226 300528 454294
rect 300208 454170 300278 454226
rect 300334 454170 300402 454226
rect 300458 454170 300528 454226
rect 300208 454102 300528 454170
rect 300208 454046 300278 454102
rect 300334 454046 300402 454102
rect 300458 454046 300528 454102
rect 300208 453978 300528 454046
rect 300208 453922 300278 453978
rect 300334 453922 300402 453978
rect 300458 453922 300528 453978
rect 300208 453888 300528 453922
rect 330928 454350 331248 454384
rect 330928 454294 330998 454350
rect 331054 454294 331122 454350
rect 331178 454294 331248 454350
rect 330928 454226 331248 454294
rect 330928 454170 330998 454226
rect 331054 454170 331122 454226
rect 331178 454170 331248 454226
rect 330928 454102 331248 454170
rect 330928 454046 330998 454102
rect 331054 454046 331122 454102
rect 331178 454046 331248 454102
rect 330928 453978 331248 454046
rect 330928 453922 330998 453978
rect 331054 453922 331122 453978
rect 331178 453922 331248 453978
rect 330928 453888 331248 453922
rect 361648 454350 361968 454384
rect 361648 454294 361718 454350
rect 361774 454294 361842 454350
rect 361898 454294 361968 454350
rect 361648 454226 361968 454294
rect 361648 454170 361718 454226
rect 361774 454170 361842 454226
rect 361898 454170 361968 454226
rect 361648 454102 361968 454170
rect 361648 454046 361718 454102
rect 361774 454046 361842 454102
rect 361898 454046 361968 454102
rect 361648 453978 361968 454046
rect 361648 453922 361718 453978
rect 361774 453922 361842 453978
rect 361898 453922 361968 453978
rect 361648 453888 361968 453922
rect 392368 454350 392688 454384
rect 392368 454294 392438 454350
rect 392494 454294 392562 454350
rect 392618 454294 392688 454350
rect 392368 454226 392688 454294
rect 392368 454170 392438 454226
rect 392494 454170 392562 454226
rect 392618 454170 392688 454226
rect 392368 454102 392688 454170
rect 392368 454046 392438 454102
rect 392494 454046 392562 454102
rect 392618 454046 392688 454102
rect 392368 453978 392688 454046
rect 392368 453922 392438 453978
rect 392494 453922 392562 453978
rect 392618 453922 392688 453978
rect 392368 453888 392688 453922
rect 423088 454350 423408 454384
rect 423088 454294 423158 454350
rect 423214 454294 423282 454350
rect 423338 454294 423408 454350
rect 423088 454226 423408 454294
rect 423088 454170 423158 454226
rect 423214 454170 423282 454226
rect 423338 454170 423408 454226
rect 423088 454102 423408 454170
rect 423088 454046 423158 454102
rect 423214 454046 423282 454102
rect 423338 454046 423408 454102
rect 423088 453978 423408 454046
rect 423088 453922 423158 453978
rect 423214 453922 423282 453978
rect 423338 453922 423408 453978
rect 423088 453888 423408 453922
rect 453808 454350 454128 454384
rect 453808 454294 453878 454350
rect 453934 454294 454002 454350
rect 454058 454294 454128 454350
rect 453808 454226 454128 454294
rect 453808 454170 453878 454226
rect 453934 454170 454002 454226
rect 454058 454170 454128 454226
rect 453808 454102 454128 454170
rect 453808 454046 453878 454102
rect 453934 454046 454002 454102
rect 454058 454046 454128 454102
rect 453808 453978 454128 454046
rect 453808 453922 453878 453978
rect 453934 453922 454002 453978
rect 454058 453922 454128 453978
rect 453808 453888 454128 453922
rect 484528 454350 484848 454384
rect 484528 454294 484598 454350
rect 484654 454294 484722 454350
rect 484778 454294 484848 454350
rect 484528 454226 484848 454294
rect 484528 454170 484598 454226
rect 484654 454170 484722 454226
rect 484778 454170 484848 454226
rect 484528 454102 484848 454170
rect 484528 454046 484598 454102
rect 484654 454046 484722 454102
rect 484778 454046 484848 454102
rect 484528 453978 484848 454046
rect 484528 453922 484598 453978
rect 484654 453922 484722 453978
rect 484778 453922 484848 453978
rect 484528 453888 484848 453922
rect 515248 454350 515568 454384
rect 515248 454294 515318 454350
rect 515374 454294 515442 454350
rect 515498 454294 515568 454350
rect 515248 454226 515568 454294
rect 515248 454170 515318 454226
rect 515374 454170 515442 454226
rect 515498 454170 515568 454226
rect 515248 454102 515568 454170
rect 515248 454046 515318 454102
rect 515374 454046 515442 454102
rect 515498 454046 515568 454102
rect 515248 453978 515568 454046
rect 515248 453922 515318 453978
rect 515374 453922 515442 453978
rect 515498 453922 515568 453978
rect 515248 453888 515568 453922
rect 545968 454350 546288 454384
rect 545968 454294 546038 454350
rect 546094 454294 546162 454350
rect 546218 454294 546288 454350
rect 545968 454226 546288 454294
rect 545968 454170 546038 454226
rect 546094 454170 546162 454226
rect 546218 454170 546288 454226
rect 545968 454102 546288 454170
rect 545968 454046 546038 454102
rect 546094 454046 546162 454102
rect 546218 454046 546288 454102
rect 545968 453978 546288 454046
rect 545968 453922 546038 453978
rect 546094 453922 546162 453978
rect 546218 453922 546288 453978
rect 545968 453888 546288 453922
rect 561154 454350 561774 471922
rect 561154 454294 561250 454350
rect 561306 454294 561374 454350
rect 561430 454294 561498 454350
rect 561554 454294 561622 454350
rect 561678 454294 561774 454350
rect 561154 454226 561774 454294
rect 561154 454170 561250 454226
rect 561306 454170 561374 454226
rect 561430 454170 561498 454226
rect 561554 454170 561622 454226
rect 561678 454170 561774 454226
rect 561154 454102 561774 454170
rect 561154 454046 561250 454102
rect 561306 454046 561374 454102
rect 561430 454046 561498 454102
rect 561554 454046 561622 454102
rect 561678 454046 561774 454102
rect 561154 453978 561774 454046
rect 561154 453922 561250 453978
rect 561306 453922 561374 453978
rect 561430 453922 561498 453978
rect 561554 453922 561622 453978
rect 561678 453922 561774 453978
rect 131248 442350 131568 442384
rect 131248 442294 131318 442350
rect 131374 442294 131442 442350
rect 131498 442294 131568 442350
rect 131248 442226 131568 442294
rect 131248 442170 131318 442226
rect 131374 442170 131442 442226
rect 131498 442170 131568 442226
rect 131248 442102 131568 442170
rect 131248 442046 131318 442102
rect 131374 442046 131442 442102
rect 131498 442046 131568 442102
rect 131248 441978 131568 442046
rect 131248 441922 131318 441978
rect 131374 441922 131442 441978
rect 131498 441922 131568 441978
rect 131248 441888 131568 441922
rect 161968 442350 162288 442384
rect 161968 442294 162038 442350
rect 162094 442294 162162 442350
rect 162218 442294 162288 442350
rect 161968 442226 162288 442294
rect 161968 442170 162038 442226
rect 162094 442170 162162 442226
rect 162218 442170 162288 442226
rect 161968 442102 162288 442170
rect 161968 442046 162038 442102
rect 162094 442046 162162 442102
rect 162218 442046 162288 442102
rect 161968 441978 162288 442046
rect 161968 441922 162038 441978
rect 162094 441922 162162 441978
rect 162218 441922 162288 441978
rect 161968 441888 162288 441922
rect 192688 442350 193008 442384
rect 192688 442294 192758 442350
rect 192814 442294 192882 442350
rect 192938 442294 193008 442350
rect 192688 442226 193008 442294
rect 192688 442170 192758 442226
rect 192814 442170 192882 442226
rect 192938 442170 193008 442226
rect 192688 442102 193008 442170
rect 192688 442046 192758 442102
rect 192814 442046 192882 442102
rect 192938 442046 193008 442102
rect 192688 441978 193008 442046
rect 192688 441922 192758 441978
rect 192814 441922 192882 441978
rect 192938 441922 193008 441978
rect 192688 441888 193008 441922
rect 223408 442350 223728 442384
rect 223408 442294 223478 442350
rect 223534 442294 223602 442350
rect 223658 442294 223728 442350
rect 223408 442226 223728 442294
rect 223408 442170 223478 442226
rect 223534 442170 223602 442226
rect 223658 442170 223728 442226
rect 223408 442102 223728 442170
rect 223408 442046 223478 442102
rect 223534 442046 223602 442102
rect 223658 442046 223728 442102
rect 223408 441978 223728 442046
rect 223408 441922 223478 441978
rect 223534 441922 223602 441978
rect 223658 441922 223728 441978
rect 223408 441888 223728 441922
rect 254128 442350 254448 442384
rect 254128 442294 254198 442350
rect 254254 442294 254322 442350
rect 254378 442294 254448 442350
rect 254128 442226 254448 442294
rect 254128 442170 254198 442226
rect 254254 442170 254322 442226
rect 254378 442170 254448 442226
rect 254128 442102 254448 442170
rect 254128 442046 254198 442102
rect 254254 442046 254322 442102
rect 254378 442046 254448 442102
rect 254128 441978 254448 442046
rect 254128 441922 254198 441978
rect 254254 441922 254322 441978
rect 254378 441922 254448 441978
rect 254128 441888 254448 441922
rect 284848 442350 285168 442384
rect 284848 442294 284918 442350
rect 284974 442294 285042 442350
rect 285098 442294 285168 442350
rect 284848 442226 285168 442294
rect 284848 442170 284918 442226
rect 284974 442170 285042 442226
rect 285098 442170 285168 442226
rect 284848 442102 285168 442170
rect 284848 442046 284918 442102
rect 284974 442046 285042 442102
rect 285098 442046 285168 442102
rect 284848 441978 285168 442046
rect 284848 441922 284918 441978
rect 284974 441922 285042 441978
rect 285098 441922 285168 441978
rect 284848 441888 285168 441922
rect 315568 442350 315888 442384
rect 315568 442294 315638 442350
rect 315694 442294 315762 442350
rect 315818 442294 315888 442350
rect 315568 442226 315888 442294
rect 315568 442170 315638 442226
rect 315694 442170 315762 442226
rect 315818 442170 315888 442226
rect 315568 442102 315888 442170
rect 315568 442046 315638 442102
rect 315694 442046 315762 442102
rect 315818 442046 315888 442102
rect 315568 441978 315888 442046
rect 315568 441922 315638 441978
rect 315694 441922 315762 441978
rect 315818 441922 315888 441978
rect 315568 441888 315888 441922
rect 346288 442350 346608 442384
rect 346288 442294 346358 442350
rect 346414 442294 346482 442350
rect 346538 442294 346608 442350
rect 346288 442226 346608 442294
rect 346288 442170 346358 442226
rect 346414 442170 346482 442226
rect 346538 442170 346608 442226
rect 346288 442102 346608 442170
rect 346288 442046 346358 442102
rect 346414 442046 346482 442102
rect 346538 442046 346608 442102
rect 346288 441978 346608 442046
rect 346288 441922 346358 441978
rect 346414 441922 346482 441978
rect 346538 441922 346608 441978
rect 346288 441888 346608 441922
rect 377008 442350 377328 442384
rect 377008 442294 377078 442350
rect 377134 442294 377202 442350
rect 377258 442294 377328 442350
rect 377008 442226 377328 442294
rect 377008 442170 377078 442226
rect 377134 442170 377202 442226
rect 377258 442170 377328 442226
rect 377008 442102 377328 442170
rect 377008 442046 377078 442102
rect 377134 442046 377202 442102
rect 377258 442046 377328 442102
rect 377008 441978 377328 442046
rect 377008 441922 377078 441978
rect 377134 441922 377202 441978
rect 377258 441922 377328 441978
rect 377008 441888 377328 441922
rect 407728 442350 408048 442384
rect 407728 442294 407798 442350
rect 407854 442294 407922 442350
rect 407978 442294 408048 442350
rect 407728 442226 408048 442294
rect 407728 442170 407798 442226
rect 407854 442170 407922 442226
rect 407978 442170 408048 442226
rect 407728 442102 408048 442170
rect 407728 442046 407798 442102
rect 407854 442046 407922 442102
rect 407978 442046 408048 442102
rect 407728 441978 408048 442046
rect 407728 441922 407798 441978
rect 407854 441922 407922 441978
rect 407978 441922 408048 441978
rect 407728 441888 408048 441922
rect 438448 442350 438768 442384
rect 438448 442294 438518 442350
rect 438574 442294 438642 442350
rect 438698 442294 438768 442350
rect 438448 442226 438768 442294
rect 438448 442170 438518 442226
rect 438574 442170 438642 442226
rect 438698 442170 438768 442226
rect 438448 442102 438768 442170
rect 438448 442046 438518 442102
rect 438574 442046 438642 442102
rect 438698 442046 438768 442102
rect 438448 441978 438768 442046
rect 438448 441922 438518 441978
rect 438574 441922 438642 441978
rect 438698 441922 438768 441978
rect 438448 441888 438768 441922
rect 469168 442350 469488 442384
rect 469168 442294 469238 442350
rect 469294 442294 469362 442350
rect 469418 442294 469488 442350
rect 469168 442226 469488 442294
rect 469168 442170 469238 442226
rect 469294 442170 469362 442226
rect 469418 442170 469488 442226
rect 469168 442102 469488 442170
rect 469168 442046 469238 442102
rect 469294 442046 469362 442102
rect 469418 442046 469488 442102
rect 469168 441978 469488 442046
rect 469168 441922 469238 441978
rect 469294 441922 469362 441978
rect 469418 441922 469488 441978
rect 469168 441888 469488 441922
rect 499888 442350 500208 442384
rect 499888 442294 499958 442350
rect 500014 442294 500082 442350
rect 500138 442294 500208 442350
rect 499888 442226 500208 442294
rect 499888 442170 499958 442226
rect 500014 442170 500082 442226
rect 500138 442170 500208 442226
rect 499888 442102 500208 442170
rect 499888 442046 499958 442102
rect 500014 442046 500082 442102
rect 500138 442046 500208 442102
rect 499888 441978 500208 442046
rect 499888 441922 499958 441978
rect 500014 441922 500082 441978
rect 500138 441922 500208 441978
rect 499888 441888 500208 441922
rect 530608 442350 530928 442384
rect 530608 442294 530678 442350
rect 530734 442294 530802 442350
rect 530858 442294 530928 442350
rect 530608 442226 530928 442294
rect 530608 442170 530678 442226
rect 530734 442170 530802 442226
rect 530858 442170 530928 442226
rect 530608 442102 530928 442170
rect 530608 442046 530678 442102
rect 530734 442046 530802 442102
rect 530858 442046 530928 442102
rect 530608 441978 530928 442046
rect 530608 441922 530678 441978
rect 530734 441922 530802 441978
rect 530858 441922 530928 441978
rect 530608 441888 530928 441922
rect 111154 436294 111250 436350
rect 111306 436294 111374 436350
rect 111430 436294 111498 436350
rect 111554 436294 111622 436350
rect 111678 436294 111774 436350
rect 111154 436226 111774 436294
rect 111154 436170 111250 436226
rect 111306 436170 111374 436226
rect 111430 436170 111498 436226
rect 111554 436170 111622 436226
rect 111678 436170 111774 436226
rect 111154 436102 111774 436170
rect 111154 436046 111250 436102
rect 111306 436046 111374 436102
rect 111430 436046 111498 436102
rect 111554 436046 111622 436102
rect 111678 436046 111774 436102
rect 111154 435978 111774 436046
rect 111154 435922 111250 435978
rect 111306 435922 111374 435978
rect 111430 435922 111498 435978
rect 111554 435922 111622 435978
rect 111678 435922 111774 435978
rect 96874 424294 96970 424350
rect 97026 424294 97094 424350
rect 97150 424294 97218 424350
rect 97274 424294 97342 424350
rect 97398 424294 97494 424350
rect 96874 424226 97494 424294
rect 96874 424170 96970 424226
rect 97026 424170 97094 424226
rect 97150 424170 97218 424226
rect 97274 424170 97342 424226
rect 97398 424170 97494 424226
rect 96874 424102 97494 424170
rect 96874 424046 96970 424102
rect 97026 424046 97094 424102
rect 97150 424046 97218 424102
rect 97274 424046 97342 424102
rect 97398 424046 97494 424102
rect 96874 423978 97494 424046
rect 96874 423922 96970 423978
rect 97026 423922 97094 423978
rect 97150 423922 97218 423978
rect 97274 423922 97342 423978
rect 97398 423922 97494 423978
rect 96874 406350 97494 423922
rect 100528 424350 100848 424384
rect 100528 424294 100598 424350
rect 100654 424294 100722 424350
rect 100778 424294 100848 424350
rect 100528 424226 100848 424294
rect 100528 424170 100598 424226
rect 100654 424170 100722 424226
rect 100778 424170 100848 424226
rect 100528 424102 100848 424170
rect 100528 424046 100598 424102
rect 100654 424046 100722 424102
rect 100778 424046 100848 424102
rect 100528 423978 100848 424046
rect 100528 423922 100598 423978
rect 100654 423922 100722 423978
rect 100778 423922 100848 423978
rect 100528 423888 100848 423922
rect 111154 418350 111774 435922
rect 115888 436350 116208 436384
rect 115888 436294 115958 436350
rect 116014 436294 116082 436350
rect 116138 436294 116208 436350
rect 115888 436226 116208 436294
rect 115888 436170 115958 436226
rect 116014 436170 116082 436226
rect 116138 436170 116208 436226
rect 115888 436102 116208 436170
rect 115888 436046 115958 436102
rect 116014 436046 116082 436102
rect 116138 436046 116208 436102
rect 115888 435978 116208 436046
rect 115888 435922 115958 435978
rect 116014 435922 116082 435978
rect 116138 435922 116208 435978
rect 115888 435888 116208 435922
rect 146608 436350 146928 436384
rect 146608 436294 146678 436350
rect 146734 436294 146802 436350
rect 146858 436294 146928 436350
rect 146608 436226 146928 436294
rect 146608 436170 146678 436226
rect 146734 436170 146802 436226
rect 146858 436170 146928 436226
rect 146608 436102 146928 436170
rect 146608 436046 146678 436102
rect 146734 436046 146802 436102
rect 146858 436046 146928 436102
rect 146608 435978 146928 436046
rect 146608 435922 146678 435978
rect 146734 435922 146802 435978
rect 146858 435922 146928 435978
rect 146608 435888 146928 435922
rect 177328 436350 177648 436384
rect 177328 436294 177398 436350
rect 177454 436294 177522 436350
rect 177578 436294 177648 436350
rect 177328 436226 177648 436294
rect 177328 436170 177398 436226
rect 177454 436170 177522 436226
rect 177578 436170 177648 436226
rect 177328 436102 177648 436170
rect 177328 436046 177398 436102
rect 177454 436046 177522 436102
rect 177578 436046 177648 436102
rect 177328 435978 177648 436046
rect 177328 435922 177398 435978
rect 177454 435922 177522 435978
rect 177578 435922 177648 435978
rect 177328 435888 177648 435922
rect 208048 436350 208368 436384
rect 208048 436294 208118 436350
rect 208174 436294 208242 436350
rect 208298 436294 208368 436350
rect 208048 436226 208368 436294
rect 208048 436170 208118 436226
rect 208174 436170 208242 436226
rect 208298 436170 208368 436226
rect 208048 436102 208368 436170
rect 208048 436046 208118 436102
rect 208174 436046 208242 436102
rect 208298 436046 208368 436102
rect 208048 435978 208368 436046
rect 208048 435922 208118 435978
rect 208174 435922 208242 435978
rect 208298 435922 208368 435978
rect 208048 435888 208368 435922
rect 238768 436350 239088 436384
rect 238768 436294 238838 436350
rect 238894 436294 238962 436350
rect 239018 436294 239088 436350
rect 238768 436226 239088 436294
rect 238768 436170 238838 436226
rect 238894 436170 238962 436226
rect 239018 436170 239088 436226
rect 238768 436102 239088 436170
rect 238768 436046 238838 436102
rect 238894 436046 238962 436102
rect 239018 436046 239088 436102
rect 238768 435978 239088 436046
rect 238768 435922 238838 435978
rect 238894 435922 238962 435978
rect 239018 435922 239088 435978
rect 238768 435888 239088 435922
rect 269488 436350 269808 436384
rect 269488 436294 269558 436350
rect 269614 436294 269682 436350
rect 269738 436294 269808 436350
rect 269488 436226 269808 436294
rect 269488 436170 269558 436226
rect 269614 436170 269682 436226
rect 269738 436170 269808 436226
rect 269488 436102 269808 436170
rect 269488 436046 269558 436102
rect 269614 436046 269682 436102
rect 269738 436046 269808 436102
rect 269488 435978 269808 436046
rect 269488 435922 269558 435978
rect 269614 435922 269682 435978
rect 269738 435922 269808 435978
rect 269488 435888 269808 435922
rect 300208 436350 300528 436384
rect 300208 436294 300278 436350
rect 300334 436294 300402 436350
rect 300458 436294 300528 436350
rect 300208 436226 300528 436294
rect 300208 436170 300278 436226
rect 300334 436170 300402 436226
rect 300458 436170 300528 436226
rect 300208 436102 300528 436170
rect 300208 436046 300278 436102
rect 300334 436046 300402 436102
rect 300458 436046 300528 436102
rect 300208 435978 300528 436046
rect 300208 435922 300278 435978
rect 300334 435922 300402 435978
rect 300458 435922 300528 435978
rect 300208 435888 300528 435922
rect 330928 436350 331248 436384
rect 330928 436294 330998 436350
rect 331054 436294 331122 436350
rect 331178 436294 331248 436350
rect 330928 436226 331248 436294
rect 330928 436170 330998 436226
rect 331054 436170 331122 436226
rect 331178 436170 331248 436226
rect 330928 436102 331248 436170
rect 330928 436046 330998 436102
rect 331054 436046 331122 436102
rect 331178 436046 331248 436102
rect 330928 435978 331248 436046
rect 330928 435922 330998 435978
rect 331054 435922 331122 435978
rect 331178 435922 331248 435978
rect 330928 435888 331248 435922
rect 361648 436350 361968 436384
rect 361648 436294 361718 436350
rect 361774 436294 361842 436350
rect 361898 436294 361968 436350
rect 361648 436226 361968 436294
rect 361648 436170 361718 436226
rect 361774 436170 361842 436226
rect 361898 436170 361968 436226
rect 361648 436102 361968 436170
rect 361648 436046 361718 436102
rect 361774 436046 361842 436102
rect 361898 436046 361968 436102
rect 361648 435978 361968 436046
rect 361648 435922 361718 435978
rect 361774 435922 361842 435978
rect 361898 435922 361968 435978
rect 361648 435888 361968 435922
rect 392368 436350 392688 436384
rect 392368 436294 392438 436350
rect 392494 436294 392562 436350
rect 392618 436294 392688 436350
rect 392368 436226 392688 436294
rect 392368 436170 392438 436226
rect 392494 436170 392562 436226
rect 392618 436170 392688 436226
rect 392368 436102 392688 436170
rect 392368 436046 392438 436102
rect 392494 436046 392562 436102
rect 392618 436046 392688 436102
rect 392368 435978 392688 436046
rect 392368 435922 392438 435978
rect 392494 435922 392562 435978
rect 392618 435922 392688 435978
rect 392368 435888 392688 435922
rect 423088 436350 423408 436384
rect 423088 436294 423158 436350
rect 423214 436294 423282 436350
rect 423338 436294 423408 436350
rect 423088 436226 423408 436294
rect 423088 436170 423158 436226
rect 423214 436170 423282 436226
rect 423338 436170 423408 436226
rect 423088 436102 423408 436170
rect 423088 436046 423158 436102
rect 423214 436046 423282 436102
rect 423338 436046 423408 436102
rect 423088 435978 423408 436046
rect 423088 435922 423158 435978
rect 423214 435922 423282 435978
rect 423338 435922 423408 435978
rect 423088 435888 423408 435922
rect 453808 436350 454128 436384
rect 453808 436294 453878 436350
rect 453934 436294 454002 436350
rect 454058 436294 454128 436350
rect 453808 436226 454128 436294
rect 453808 436170 453878 436226
rect 453934 436170 454002 436226
rect 454058 436170 454128 436226
rect 453808 436102 454128 436170
rect 453808 436046 453878 436102
rect 453934 436046 454002 436102
rect 454058 436046 454128 436102
rect 453808 435978 454128 436046
rect 453808 435922 453878 435978
rect 453934 435922 454002 435978
rect 454058 435922 454128 435978
rect 453808 435888 454128 435922
rect 484528 436350 484848 436384
rect 484528 436294 484598 436350
rect 484654 436294 484722 436350
rect 484778 436294 484848 436350
rect 484528 436226 484848 436294
rect 484528 436170 484598 436226
rect 484654 436170 484722 436226
rect 484778 436170 484848 436226
rect 484528 436102 484848 436170
rect 484528 436046 484598 436102
rect 484654 436046 484722 436102
rect 484778 436046 484848 436102
rect 484528 435978 484848 436046
rect 484528 435922 484598 435978
rect 484654 435922 484722 435978
rect 484778 435922 484848 435978
rect 484528 435888 484848 435922
rect 515248 436350 515568 436384
rect 515248 436294 515318 436350
rect 515374 436294 515442 436350
rect 515498 436294 515568 436350
rect 515248 436226 515568 436294
rect 515248 436170 515318 436226
rect 515374 436170 515442 436226
rect 515498 436170 515568 436226
rect 515248 436102 515568 436170
rect 515248 436046 515318 436102
rect 515374 436046 515442 436102
rect 515498 436046 515568 436102
rect 515248 435978 515568 436046
rect 515248 435922 515318 435978
rect 515374 435922 515442 435978
rect 515498 435922 515568 435978
rect 515248 435888 515568 435922
rect 545968 436350 546288 436384
rect 545968 436294 546038 436350
rect 546094 436294 546162 436350
rect 546218 436294 546288 436350
rect 545968 436226 546288 436294
rect 545968 436170 546038 436226
rect 546094 436170 546162 436226
rect 546218 436170 546288 436226
rect 545968 436102 546288 436170
rect 545968 436046 546038 436102
rect 546094 436046 546162 436102
rect 546218 436046 546288 436102
rect 545968 435978 546288 436046
rect 545968 435922 546038 435978
rect 546094 435922 546162 435978
rect 546218 435922 546288 435978
rect 545968 435888 546288 435922
rect 561154 436350 561774 453922
rect 561154 436294 561250 436350
rect 561306 436294 561374 436350
rect 561430 436294 561498 436350
rect 561554 436294 561622 436350
rect 561678 436294 561774 436350
rect 561154 436226 561774 436294
rect 561154 436170 561250 436226
rect 561306 436170 561374 436226
rect 561430 436170 561498 436226
rect 561554 436170 561622 436226
rect 561678 436170 561774 436226
rect 561154 436102 561774 436170
rect 561154 436046 561250 436102
rect 561306 436046 561374 436102
rect 561430 436046 561498 436102
rect 561554 436046 561622 436102
rect 561678 436046 561774 436102
rect 561154 435978 561774 436046
rect 561154 435922 561250 435978
rect 561306 435922 561374 435978
rect 561430 435922 561498 435978
rect 561554 435922 561622 435978
rect 561678 435922 561774 435978
rect 131248 424350 131568 424384
rect 131248 424294 131318 424350
rect 131374 424294 131442 424350
rect 131498 424294 131568 424350
rect 131248 424226 131568 424294
rect 131248 424170 131318 424226
rect 131374 424170 131442 424226
rect 131498 424170 131568 424226
rect 131248 424102 131568 424170
rect 131248 424046 131318 424102
rect 131374 424046 131442 424102
rect 131498 424046 131568 424102
rect 131248 423978 131568 424046
rect 131248 423922 131318 423978
rect 131374 423922 131442 423978
rect 131498 423922 131568 423978
rect 131248 423888 131568 423922
rect 161968 424350 162288 424384
rect 161968 424294 162038 424350
rect 162094 424294 162162 424350
rect 162218 424294 162288 424350
rect 161968 424226 162288 424294
rect 161968 424170 162038 424226
rect 162094 424170 162162 424226
rect 162218 424170 162288 424226
rect 161968 424102 162288 424170
rect 161968 424046 162038 424102
rect 162094 424046 162162 424102
rect 162218 424046 162288 424102
rect 161968 423978 162288 424046
rect 161968 423922 162038 423978
rect 162094 423922 162162 423978
rect 162218 423922 162288 423978
rect 161968 423888 162288 423922
rect 192688 424350 193008 424384
rect 192688 424294 192758 424350
rect 192814 424294 192882 424350
rect 192938 424294 193008 424350
rect 192688 424226 193008 424294
rect 192688 424170 192758 424226
rect 192814 424170 192882 424226
rect 192938 424170 193008 424226
rect 192688 424102 193008 424170
rect 192688 424046 192758 424102
rect 192814 424046 192882 424102
rect 192938 424046 193008 424102
rect 192688 423978 193008 424046
rect 192688 423922 192758 423978
rect 192814 423922 192882 423978
rect 192938 423922 193008 423978
rect 192688 423888 193008 423922
rect 223408 424350 223728 424384
rect 223408 424294 223478 424350
rect 223534 424294 223602 424350
rect 223658 424294 223728 424350
rect 223408 424226 223728 424294
rect 223408 424170 223478 424226
rect 223534 424170 223602 424226
rect 223658 424170 223728 424226
rect 223408 424102 223728 424170
rect 223408 424046 223478 424102
rect 223534 424046 223602 424102
rect 223658 424046 223728 424102
rect 223408 423978 223728 424046
rect 223408 423922 223478 423978
rect 223534 423922 223602 423978
rect 223658 423922 223728 423978
rect 223408 423888 223728 423922
rect 254128 424350 254448 424384
rect 254128 424294 254198 424350
rect 254254 424294 254322 424350
rect 254378 424294 254448 424350
rect 254128 424226 254448 424294
rect 254128 424170 254198 424226
rect 254254 424170 254322 424226
rect 254378 424170 254448 424226
rect 254128 424102 254448 424170
rect 254128 424046 254198 424102
rect 254254 424046 254322 424102
rect 254378 424046 254448 424102
rect 254128 423978 254448 424046
rect 254128 423922 254198 423978
rect 254254 423922 254322 423978
rect 254378 423922 254448 423978
rect 254128 423888 254448 423922
rect 284848 424350 285168 424384
rect 284848 424294 284918 424350
rect 284974 424294 285042 424350
rect 285098 424294 285168 424350
rect 284848 424226 285168 424294
rect 284848 424170 284918 424226
rect 284974 424170 285042 424226
rect 285098 424170 285168 424226
rect 284848 424102 285168 424170
rect 284848 424046 284918 424102
rect 284974 424046 285042 424102
rect 285098 424046 285168 424102
rect 284848 423978 285168 424046
rect 284848 423922 284918 423978
rect 284974 423922 285042 423978
rect 285098 423922 285168 423978
rect 284848 423888 285168 423922
rect 315568 424350 315888 424384
rect 315568 424294 315638 424350
rect 315694 424294 315762 424350
rect 315818 424294 315888 424350
rect 315568 424226 315888 424294
rect 315568 424170 315638 424226
rect 315694 424170 315762 424226
rect 315818 424170 315888 424226
rect 315568 424102 315888 424170
rect 315568 424046 315638 424102
rect 315694 424046 315762 424102
rect 315818 424046 315888 424102
rect 315568 423978 315888 424046
rect 315568 423922 315638 423978
rect 315694 423922 315762 423978
rect 315818 423922 315888 423978
rect 315568 423888 315888 423922
rect 346288 424350 346608 424384
rect 346288 424294 346358 424350
rect 346414 424294 346482 424350
rect 346538 424294 346608 424350
rect 346288 424226 346608 424294
rect 346288 424170 346358 424226
rect 346414 424170 346482 424226
rect 346538 424170 346608 424226
rect 346288 424102 346608 424170
rect 346288 424046 346358 424102
rect 346414 424046 346482 424102
rect 346538 424046 346608 424102
rect 346288 423978 346608 424046
rect 346288 423922 346358 423978
rect 346414 423922 346482 423978
rect 346538 423922 346608 423978
rect 346288 423888 346608 423922
rect 377008 424350 377328 424384
rect 377008 424294 377078 424350
rect 377134 424294 377202 424350
rect 377258 424294 377328 424350
rect 377008 424226 377328 424294
rect 377008 424170 377078 424226
rect 377134 424170 377202 424226
rect 377258 424170 377328 424226
rect 377008 424102 377328 424170
rect 377008 424046 377078 424102
rect 377134 424046 377202 424102
rect 377258 424046 377328 424102
rect 377008 423978 377328 424046
rect 377008 423922 377078 423978
rect 377134 423922 377202 423978
rect 377258 423922 377328 423978
rect 377008 423888 377328 423922
rect 407728 424350 408048 424384
rect 407728 424294 407798 424350
rect 407854 424294 407922 424350
rect 407978 424294 408048 424350
rect 407728 424226 408048 424294
rect 407728 424170 407798 424226
rect 407854 424170 407922 424226
rect 407978 424170 408048 424226
rect 407728 424102 408048 424170
rect 407728 424046 407798 424102
rect 407854 424046 407922 424102
rect 407978 424046 408048 424102
rect 407728 423978 408048 424046
rect 407728 423922 407798 423978
rect 407854 423922 407922 423978
rect 407978 423922 408048 423978
rect 407728 423888 408048 423922
rect 438448 424350 438768 424384
rect 438448 424294 438518 424350
rect 438574 424294 438642 424350
rect 438698 424294 438768 424350
rect 438448 424226 438768 424294
rect 438448 424170 438518 424226
rect 438574 424170 438642 424226
rect 438698 424170 438768 424226
rect 438448 424102 438768 424170
rect 438448 424046 438518 424102
rect 438574 424046 438642 424102
rect 438698 424046 438768 424102
rect 438448 423978 438768 424046
rect 438448 423922 438518 423978
rect 438574 423922 438642 423978
rect 438698 423922 438768 423978
rect 438448 423888 438768 423922
rect 469168 424350 469488 424384
rect 469168 424294 469238 424350
rect 469294 424294 469362 424350
rect 469418 424294 469488 424350
rect 469168 424226 469488 424294
rect 469168 424170 469238 424226
rect 469294 424170 469362 424226
rect 469418 424170 469488 424226
rect 469168 424102 469488 424170
rect 469168 424046 469238 424102
rect 469294 424046 469362 424102
rect 469418 424046 469488 424102
rect 469168 423978 469488 424046
rect 469168 423922 469238 423978
rect 469294 423922 469362 423978
rect 469418 423922 469488 423978
rect 469168 423888 469488 423922
rect 499888 424350 500208 424384
rect 499888 424294 499958 424350
rect 500014 424294 500082 424350
rect 500138 424294 500208 424350
rect 499888 424226 500208 424294
rect 499888 424170 499958 424226
rect 500014 424170 500082 424226
rect 500138 424170 500208 424226
rect 499888 424102 500208 424170
rect 499888 424046 499958 424102
rect 500014 424046 500082 424102
rect 500138 424046 500208 424102
rect 499888 423978 500208 424046
rect 499888 423922 499958 423978
rect 500014 423922 500082 423978
rect 500138 423922 500208 423978
rect 499888 423888 500208 423922
rect 530608 424350 530928 424384
rect 530608 424294 530678 424350
rect 530734 424294 530802 424350
rect 530858 424294 530928 424350
rect 530608 424226 530928 424294
rect 530608 424170 530678 424226
rect 530734 424170 530802 424226
rect 530858 424170 530928 424226
rect 530608 424102 530928 424170
rect 530608 424046 530678 424102
rect 530734 424046 530802 424102
rect 530858 424046 530928 424102
rect 530608 423978 530928 424046
rect 530608 423922 530678 423978
rect 530734 423922 530802 423978
rect 530858 423922 530928 423978
rect 530608 423888 530928 423922
rect 111154 418294 111250 418350
rect 111306 418294 111374 418350
rect 111430 418294 111498 418350
rect 111554 418294 111622 418350
rect 111678 418294 111774 418350
rect 111154 418226 111774 418294
rect 111154 418170 111250 418226
rect 111306 418170 111374 418226
rect 111430 418170 111498 418226
rect 111554 418170 111622 418226
rect 111678 418170 111774 418226
rect 111154 418102 111774 418170
rect 111154 418046 111250 418102
rect 111306 418046 111374 418102
rect 111430 418046 111498 418102
rect 111554 418046 111622 418102
rect 111678 418046 111774 418102
rect 111154 417978 111774 418046
rect 111154 417922 111250 417978
rect 111306 417922 111374 417978
rect 111430 417922 111498 417978
rect 111554 417922 111622 417978
rect 111678 417922 111774 417978
rect 96874 406294 96970 406350
rect 97026 406294 97094 406350
rect 97150 406294 97218 406350
rect 97274 406294 97342 406350
rect 97398 406294 97494 406350
rect 96874 406226 97494 406294
rect 96874 406170 96970 406226
rect 97026 406170 97094 406226
rect 97150 406170 97218 406226
rect 97274 406170 97342 406226
rect 97398 406170 97494 406226
rect 96874 406102 97494 406170
rect 96874 406046 96970 406102
rect 97026 406046 97094 406102
rect 97150 406046 97218 406102
rect 97274 406046 97342 406102
rect 97398 406046 97494 406102
rect 96874 405978 97494 406046
rect 96874 405922 96970 405978
rect 97026 405922 97094 405978
rect 97150 405922 97218 405978
rect 97274 405922 97342 405978
rect 97398 405922 97494 405978
rect 96874 388350 97494 405922
rect 100528 406350 100848 406384
rect 100528 406294 100598 406350
rect 100654 406294 100722 406350
rect 100778 406294 100848 406350
rect 100528 406226 100848 406294
rect 100528 406170 100598 406226
rect 100654 406170 100722 406226
rect 100778 406170 100848 406226
rect 100528 406102 100848 406170
rect 100528 406046 100598 406102
rect 100654 406046 100722 406102
rect 100778 406046 100848 406102
rect 100528 405978 100848 406046
rect 100528 405922 100598 405978
rect 100654 405922 100722 405978
rect 100778 405922 100848 405978
rect 100528 405888 100848 405922
rect 111154 400350 111774 417922
rect 115888 418350 116208 418384
rect 115888 418294 115958 418350
rect 116014 418294 116082 418350
rect 116138 418294 116208 418350
rect 115888 418226 116208 418294
rect 115888 418170 115958 418226
rect 116014 418170 116082 418226
rect 116138 418170 116208 418226
rect 115888 418102 116208 418170
rect 115888 418046 115958 418102
rect 116014 418046 116082 418102
rect 116138 418046 116208 418102
rect 115888 417978 116208 418046
rect 115888 417922 115958 417978
rect 116014 417922 116082 417978
rect 116138 417922 116208 417978
rect 115888 417888 116208 417922
rect 146608 418350 146928 418384
rect 146608 418294 146678 418350
rect 146734 418294 146802 418350
rect 146858 418294 146928 418350
rect 146608 418226 146928 418294
rect 146608 418170 146678 418226
rect 146734 418170 146802 418226
rect 146858 418170 146928 418226
rect 146608 418102 146928 418170
rect 146608 418046 146678 418102
rect 146734 418046 146802 418102
rect 146858 418046 146928 418102
rect 146608 417978 146928 418046
rect 146608 417922 146678 417978
rect 146734 417922 146802 417978
rect 146858 417922 146928 417978
rect 146608 417888 146928 417922
rect 177328 418350 177648 418384
rect 177328 418294 177398 418350
rect 177454 418294 177522 418350
rect 177578 418294 177648 418350
rect 177328 418226 177648 418294
rect 177328 418170 177398 418226
rect 177454 418170 177522 418226
rect 177578 418170 177648 418226
rect 177328 418102 177648 418170
rect 177328 418046 177398 418102
rect 177454 418046 177522 418102
rect 177578 418046 177648 418102
rect 177328 417978 177648 418046
rect 177328 417922 177398 417978
rect 177454 417922 177522 417978
rect 177578 417922 177648 417978
rect 177328 417888 177648 417922
rect 208048 418350 208368 418384
rect 208048 418294 208118 418350
rect 208174 418294 208242 418350
rect 208298 418294 208368 418350
rect 208048 418226 208368 418294
rect 208048 418170 208118 418226
rect 208174 418170 208242 418226
rect 208298 418170 208368 418226
rect 208048 418102 208368 418170
rect 208048 418046 208118 418102
rect 208174 418046 208242 418102
rect 208298 418046 208368 418102
rect 208048 417978 208368 418046
rect 208048 417922 208118 417978
rect 208174 417922 208242 417978
rect 208298 417922 208368 417978
rect 208048 417888 208368 417922
rect 238768 418350 239088 418384
rect 238768 418294 238838 418350
rect 238894 418294 238962 418350
rect 239018 418294 239088 418350
rect 238768 418226 239088 418294
rect 238768 418170 238838 418226
rect 238894 418170 238962 418226
rect 239018 418170 239088 418226
rect 238768 418102 239088 418170
rect 238768 418046 238838 418102
rect 238894 418046 238962 418102
rect 239018 418046 239088 418102
rect 238768 417978 239088 418046
rect 238768 417922 238838 417978
rect 238894 417922 238962 417978
rect 239018 417922 239088 417978
rect 238768 417888 239088 417922
rect 269488 418350 269808 418384
rect 269488 418294 269558 418350
rect 269614 418294 269682 418350
rect 269738 418294 269808 418350
rect 269488 418226 269808 418294
rect 269488 418170 269558 418226
rect 269614 418170 269682 418226
rect 269738 418170 269808 418226
rect 269488 418102 269808 418170
rect 269488 418046 269558 418102
rect 269614 418046 269682 418102
rect 269738 418046 269808 418102
rect 269488 417978 269808 418046
rect 269488 417922 269558 417978
rect 269614 417922 269682 417978
rect 269738 417922 269808 417978
rect 269488 417888 269808 417922
rect 300208 418350 300528 418384
rect 300208 418294 300278 418350
rect 300334 418294 300402 418350
rect 300458 418294 300528 418350
rect 300208 418226 300528 418294
rect 300208 418170 300278 418226
rect 300334 418170 300402 418226
rect 300458 418170 300528 418226
rect 300208 418102 300528 418170
rect 300208 418046 300278 418102
rect 300334 418046 300402 418102
rect 300458 418046 300528 418102
rect 300208 417978 300528 418046
rect 300208 417922 300278 417978
rect 300334 417922 300402 417978
rect 300458 417922 300528 417978
rect 300208 417888 300528 417922
rect 330928 418350 331248 418384
rect 330928 418294 330998 418350
rect 331054 418294 331122 418350
rect 331178 418294 331248 418350
rect 330928 418226 331248 418294
rect 330928 418170 330998 418226
rect 331054 418170 331122 418226
rect 331178 418170 331248 418226
rect 330928 418102 331248 418170
rect 330928 418046 330998 418102
rect 331054 418046 331122 418102
rect 331178 418046 331248 418102
rect 330928 417978 331248 418046
rect 330928 417922 330998 417978
rect 331054 417922 331122 417978
rect 331178 417922 331248 417978
rect 330928 417888 331248 417922
rect 361648 418350 361968 418384
rect 361648 418294 361718 418350
rect 361774 418294 361842 418350
rect 361898 418294 361968 418350
rect 361648 418226 361968 418294
rect 361648 418170 361718 418226
rect 361774 418170 361842 418226
rect 361898 418170 361968 418226
rect 361648 418102 361968 418170
rect 361648 418046 361718 418102
rect 361774 418046 361842 418102
rect 361898 418046 361968 418102
rect 361648 417978 361968 418046
rect 361648 417922 361718 417978
rect 361774 417922 361842 417978
rect 361898 417922 361968 417978
rect 361648 417888 361968 417922
rect 392368 418350 392688 418384
rect 392368 418294 392438 418350
rect 392494 418294 392562 418350
rect 392618 418294 392688 418350
rect 392368 418226 392688 418294
rect 392368 418170 392438 418226
rect 392494 418170 392562 418226
rect 392618 418170 392688 418226
rect 392368 418102 392688 418170
rect 392368 418046 392438 418102
rect 392494 418046 392562 418102
rect 392618 418046 392688 418102
rect 392368 417978 392688 418046
rect 392368 417922 392438 417978
rect 392494 417922 392562 417978
rect 392618 417922 392688 417978
rect 392368 417888 392688 417922
rect 423088 418350 423408 418384
rect 423088 418294 423158 418350
rect 423214 418294 423282 418350
rect 423338 418294 423408 418350
rect 423088 418226 423408 418294
rect 423088 418170 423158 418226
rect 423214 418170 423282 418226
rect 423338 418170 423408 418226
rect 423088 418102 423408 418170
rect 423088 418046 423158 418102
rect 423214 418046 423282 418102
rect 423338 418046 423408 418102
rect 423088 417978 423408 418046
rect 423088 417922 423158 417978
rect 423214 417922 423282 417978
rect 423338 417922 423408 417978
rect 423088 417888 423408 417922
rect 453808 418350 454128 418384
rect 453808 418294 453878 418350
rect 453934 418294 454002 418350
rect 454058 418294 454128 418350
rect 453808 418226 454128 418294
rect 453808 418170 453878 418226
rect 453934 418170 454002 418226
rect 454058 418170 454128 418226
rect 453808 418102 454128 418170
rect 453808 418046 453878 418102
rect 453934 418046 454002 418102
rect 454058 418046 454128 418102
rect 453808 417978 454128 418046
rect 453808 417922 453878 417978
rect 453934 417922 454002 417978
rect 454058 417922 454128 417978
rect 453808 417888 454128 417922
rect 484528 418350 484848 418384
rect 484528 418294 484598 418350
rect 484654 418294 484722 418350
rect 484778 418294 484848 418350
rect 484528 418226 484848 418294
rect 484528 418170 484598 418226
rect 484654 418170 484722 418226
rect 484778 418170 484848 418226
rect 484528 418102 484848 418170
rect 484528 418046 484598 418102
rect 484654 418046 484722 418102
rect 484778 418046 484848 418102
rect 484528 417978 484848 418046
rect 484528 417922 484598 417978
rect 484654 417922 484722 417978
rect 484778 417922 484848 417978
rect 484528 417888 484848 417922
rect 515248 418350 515568 418384
rect 515248 418294 515318 418350
rect 515374 418294 515442 418350
rect 515498 418294 515568 418350
rect 515248 418226 515568 418294
rect 515248 418170 515318 418226
rect 515374 418170 515442 418226
rect 515498 418170 515568 418226
rect 515248 418102 515568 418170
rect 515248 418046 515318 418102
rect 515374 418046 515442 418102
rect 515498 418046 515568 418102
rect 515248 417978 515568 418046
rect 515248 417922 515318 417978
rect 515374 417922 515442 417978
rect 515498 417922 515568 417978
rect 515248 417888 515568 417922
rect 545968 418350 546288 418384
rect 545968 418294 546038 418350
rect 546094 418294 546162 418350
rect 546218 418294 546288 418350
rect 545968 418226 546288 418294
rect 545968 418170 546038 418226
rect 546094 418170 546162 418226
rect 546218 418170 546288 418226
rect 545968 418102 546288 418170
rect 545968 418046 546038 418102
rect 546094 418046 546162 418102
rect 546218 418046 546288 418102
rect 545968 417978 546288 418046
rect 545968 417922 546038 417978
rect 546094 417922 546162 417978
rect 546218 417922 546288 417978
rect 545968 417888 546288 417922
rect 561154 418350 561774 435922
rect 561154 418294 561250 418350
rect 561306 418294 561374 418350
rect 561430 418294 561498 418350
rect 561554 418294 561622 418350
rect 561678 418294 561774 418350
rect 561154 418226 561774 418294
rect 561154 418170 561250 418226
rect 561306 418170 561374 418226
rect 561430 418170 561498 418226
rect 561554 418170 561622 418226
rect 561678 418170 561774 418226
rect 561154 418102 561774 418170
rect 561154 418046 561250 418102
rect 561306 418046 561374 418102
rect 561430 418046 561498 418102
rect 561554 418046 561622 418102
rect 561678 418046 561774 418102
rect 561154 417978 561774 418046
rect 561154 417922 561250 417978
rect 561306 417922 561374 417978
rect 561430 417922 561498 417978
rect 561554 417922 561622 417978
rect 561678 417922 561774 417978
rect 131248 406350 131568 406384
rect 131248 406294 131318 406350
rect 131374 406294 131442 406350
rect 131498 406294 131568 406350
rect 131248 406226 131568 406294
rect 131248 406170 131318 406226
rect 131374 406170 131442 406226
rect 131498 406170 131568 406226
rect 131248 406102 131568 406170
rect 131248 406046 131318 406102
rect 131374 406046 131442 406102
rect 131498 406046 131568 406102
rect 131248 405978 131568 406046
rect 131248 405922 131318 405978
rect 131374 405922 131442 405978
rect 131498 405922 131568 405978
rect 131248 405888 131568 405922
rect 161968 406350 162288 406384
rect 161968 406294 162038 406350
rect 162094 406294 162162 406350
rect 162218 406294 162288 406350
rect 161968 406226 162288 406294
rect 161968 406170 162038 406226
rect 162094 406170 162162 406226
rect 162218 406170 162288 406226
rect 161968 406102 162288 406170
rect 161968 406046 162038 406102
rect 162094 406046 162162 406102
rect 162218 406046 162288 406102
rect 161968 405978 162288 406046
rect 161968 405922 162038 405978
rect 162094 405922 162162 405978
rect 162218 405922 162288 405978
rect 161968 405888 162288 405922
rect 192688 406350 193008 406384
rect 192688 406294 192758 406350
rect 192814 406294 192882 406350
rect 192938 406294 193008 406350
rect 192688 406226 193008 406294
rect 192688 406170 192758 406226
rect 192814 406170 192882 406226
rect 192938 406170 193008 406226
rect 192688 406102 193008 406170
rect 192688 406046 192758 406102
rect 192814 406046 192882 406102
rect 192938 406046 193008 406102
rect 192688 405978 193008 406046
rect 192688 405922 192758 405978
rect 192814 405922 192882 405978
rect 192938 405922 193008 405978
rect 192688 405888 193008 405922
rect 223408 406350 223728 406384
rect 223408 406294 223478 406350
rect 223534 406294 223602 406350
rect 223658 406294 223728 406350
rect 223408 406226 223728 406294
rect 223408 406170 223478 406226
rect 223534 406170 223602 406226
rect 223658 406170 223728 406226
rect 223408 406102 223728 406170
rect 223408 406046 223478 406102
rect 223534 406046 223602 406102
rect 223658 406046 223728 406102
rect 223408 405978 223728 406046
rect 223408 405922 223478 405978
rect 223534 405922 223602 405978
rect 223658 405922 223728 405978
rect 223408 405888 223728 405922
rect 254128 406350 254448 406384
rect 254128 406294 254198 406350
rect 254254 406294 254322 406350
rect 254378 406294 254448 406350
rect 254128 406226 254448 406294
rect 254128 406170 254198 406226
rect 254254 406170 254322 406226
rect 254378 406170 254448 406226
rect 254128 406102 254448 406170
rect 254128 406046 254198 406102
rect 254254 406046 254322 406102
rect 254378 406046 254448 406102
rect 254128 405978 254448 406046
rect 254128 405922 254198 405978
rect 254254 405922 254322 405978
rect 254378 405922 254448 405978
rect 254128 405888 254448 405922
rect 284848 406350 285168 406384
rect 284848 406294 284918 406350
rect 284974 406294 285042 406350
rect 285098 406294 285168 406350
rect 284848 406226 285168 406294
rect 284848 406170 284918 406226
rect 284974 406170 285042 406226
rect 285098 406170 285168 406226
rect 284848 406102 285168 406170
rect 284848 406046 284918 406102
rect 284974 406046 285042 406102
rect 285098 406046 285168 406102
rect 284848 405978 285168 406046
rect 284848 405922 284918 405978
rect 284974 405922 285042 405978
rect 285098 405922 285168 405978
rect 284848 405888 285168 405922
rect 315568 406350 315888 406384
rect 315568 406294 315638 406350
rect 315694 406294 315762 406350
rect 315818 406294 315888 406350
rect 315568 406226 315888 406294
rect 315568 406170 315638 406226
rect 315694 406170 315762 406226
rect 315818 406170 315888 406226
rect 315568 406102 315888 406170
rect 315568 406046 315638 406102
rect 315694 406046 315762 406102
rect 315818 406046 315888 406102
rect 315568 405978 315888 406046
rect 315568 405922 315638 405978
rect 315694 405922 315762 405978
rect 315818 405922 315888 405978
rect 315568 405888 315888 405922
rect 346288 406350 346608 406384
rect 346288 406294 346358 406350
rect 346414 406294 346482 406350
rect 346538 406294 346608 406350
rect 346288 406226 346608 406294
rect 346288 406170 346358 406226
rect 346414 406170 346482 406226
rect 346538 406170 346608 406226
rect 346288 406102 346608 406170
rect 346288 406046 346358 406102
rect 346414 406046 346482 406102
rect 346538 406046 346608 406102
rect 346288 405978 346608 406046
rect 346288 405922 346358 405978
rect 346414 405922 346482 405978
rect 346538 405922 346608 405978
rect 346288 405888 346608 405922
rect 377008 406350 377328 406384
rect 377008 406294 377078 406350
rect 377134 406294 377202 406350
rect 377258 406294 377328 406350
rect 377008 406226 377328 406294
rect 377008 406170 377078 406226
rect 377134 406170 377202 406226
rect 377258 406170 377328 406226
rect 377008 406102 377328 406170
rect 377008 406046 377078 406102
rect 377134 406046 377202 406102
rect 377258 406046 377328 406102
rect 377008 405978 377328 406046
rect 377008 405922 377078 405978
rect 377134 405922 377202 405978
rect 377258 405922 377328 405978
rect 377008 405888 377328 405922
rect 407728 406350 408048 406384
rect 407728 406294 407798 406350
rect 407854 406294 407922 406350
rect 407978 406294 408048 406350
rect 407728 406226 408048 406294
rect 407728 406170 407798 406226
rect 407854 406170 407922 406226
rect 407978 406170 408048 406226
rect 407728 406102 408048 406170
rect 407728 406046 407798 406102
rect 407854 406046 407922 406102
rect 407978 406046 408048 406102
rect 407728 405978 408048 406046
rect 407728 405922 407798 405978
rect 407854 405922 407922 405978
rect 407978 405922 408048 405978
rect 407728 405888 408048 405922
rect 438448 406350 438768 406384
rect 438448 406294 438518 406350
rect 438574 406294 438642 406350
rect 438698 406294 438768 406350
rect 438448 406226 438768 406294
rect 438448 406170 438518 406226
rect 438574 406170 438642 406226
rect 438698 406170 438768 406226
rect 438448 406102 438768 406170
rect 438448 406046 438518 406102
rect 438574 406046 438642 406102
rect 438698 406046 438768 406102
rect 438448 405978 438768 406046
rect 438448 405922 438518 405978
rect 438574 405922 438642 405978
rect 438698 405922 438768 405978
rect 438448 405888 438768 405922
rect 469168 406350 469488 406384
rect 469168 406294 469238 406350
rect 469294 406294 469362 406350
rect 469418 406294 469488 406350
rect 469168 406226 469488 406294
rect 469168 406170 469238 406226
rect 469294 406170 469362 406226
rect 469418 406170 469488 406226
rect 469168 406102 469488 406170
rect 469168 406046 469238 406102
rect 469294 406046 469362 406102
rect 469418 406046 469488 406102
rect 469168 405978 469488 406046
rect 469168 405922 469238 405978
rect 469294 405922 469362 405978
rect 469418 405922 469488 405978
rect 469168 405888 469488 405922
rect 499888 406350 500208 406384
rect 499888 406294 499958 406350
rect 500014 406294 500082 406350
rect 500138 406294 500208 406350
rect 499888 406226 500208 406294
rect 499888 406170 499958 406226
rect 500014 406170 500082 406226
rect 500138 406170 500208 406226
rect 499888 406102 500208 406170
rect 499888 406046 499958 406102
rect 500014 406046 500082 406102
rect 500138 406046 500208 406102
rect 499888 405978 500208 406046
rect 499888 405922 499958 405978
rect 500014 405922 500082 405978
rect 500138 405922 500208 405978
rect 499888 405888 500208 405922
rect 530608 406350 530928 406384
rect 530608 406294 530678 406350
rect 530734 406294 530802 406350
rect 530858 406294 530928 406350
rect 530608 406226 530928 406294
rect 530608 406170 530678 406226
rect 530734 406170 530802 406226
rect 530858 406170 530928 406226
rect 530608 406102 530928 406170
rect 530608 406046 530678 406102
rect 530734 406046 530802 406102
rect 530858 406046 530928 406102
rect 530608 405978 530928 406046
rect 530608 405922 530678 405978
rect 530734 405922 530802 405978
rect 530858 405922 530928 405978
rect 530608 405888 530928 405922
rect 111154 400294 111250 400350
rect 111306 400294 111374 400350
rect 111430 400294 111498 400350
rect 111554 400294 111622 400350
rect 111678 400294 111774 400350
rect 111154 400226 111774 400294
rect 111154 400170 111250 400226
rect 111306 400170 111374 400226
rect 111430 400170 111498 400226
rect 111554 400170 111622 400226
rect 111678 400170 111774 400226
rect 111154 400102 111774 400170
rect 111154 400046 111250 400102
rect 111306 400046 111374 400102
rect 111430 400046 111498 400102
rect 111554 400046 111622 400102
rect 111678 400046 111774 400102
rect 111154 399978 111774 400046
rect 111154 399922 111250 399978
rect 111306 399922 111374 399978
rect 111430 399922 111498 399978
rect 111554 399922 111622 399978
rect 111678 399922 111774 399978
rect 96874 388294 96970 388350
rect 97026 388294 97094 388350
rect 97150 388294 97218 388350
rect 97274 388294 97342 388350
rect 97398 388294 97494 388350
rect 96874 388226 97494 388294
rect 96874 388170 96970 388226
rect 97026 388170 97094 388226
rect 97150 388170 97218 388226
rect 97274 388170 97342 388226
rect 97398 388170 97494 388226
rect 96874 388102 97494 388170
rect 96874 388046 96970 388102
rect 97026 388046 97094 388102
rect 97150 388046 97218 388102
rect 97274 388046 97342 388102
rect 97398 388046 97494 388102
rect 96874 387978 97494 388046
rect 96874 387922 96970 387978
rect 97026 387922 97094 387978
rect 97150 387922 97218 387978
rect 97274 387922 97342 387978
rect 97398 387922 97494 387978
rect 96874 370350 97494 387922
rect 100528 388350 100848 388384
rect 100528 388294 100598 388350
rect 100654 388294 100722 388350
rect 100778 388294 100848 388350
rect 100528 388226 100848 388294
rect 100528 388170 100598 388226
rect 100654 388170 100722 388226
rect 100778 388170 100848 388226
rect 100528 388102 100848 388170
rect 100528 388046 100598 388102
rect 100654 388046 100722 388102
rect 100778 388046 100848 388102
rect 100528 387978 100848 388046
rect 100528 387922 100598 387978
rect 100654 387922 100722 387978
rect 100778 387922 100848 387978
rect 100528 387888 100848 387922
rect 111154 382350 111774 399922
rect 115888 400350 116208 400384
rect 115888 400294 115958 400350
rect 116014 400294 116082 400350
rect 116138 400294 116208 400350
rect 115888 400226 116208 400294
rect 115888 400170 115958 400226
rect 116014 400170 116082 400226
rect 116138 400170 116208 400226
rect 115888 400102 116208 400170
rect 115888 400046 115958 400102
rect 116014 400046 116082 400102
rect 116138 400046 116208 400102
rect 115888 399978 116208 400046
rect 115888 399922 115958 399978
rect 116014 399922 116082 399978
rect 116138 399922 116208 399978
rect 115888 399888 116208 399922
rect 146608 400350 146928 400384
rect 146608 400294 146678 400350
rect 146734 400294 146802 400350
rect 146858 400294 146928 400350
rect 146608 400226 146928 400294
rect 146608 400170 146678 400226
rect 146734 400170 146802 400226
rect 146858 400170 146928 400226
rect 146608 400102 146928 400170
rect 146608 400046 146678 400102
rect 146734 400046 146802 400102
rect 146858 400046 146928 400102
rect 146608 399978 146928 400046
rect 146608 399922 146678 399978
rect 146734 399922 146802 399978
rect 146858 399922 146928 399978
rect 146608 399888 146928 399922
rect 177328 400350 177648 400384
rect 177328 400294 177398 400350
rect 177454 400294 177522 400350
rect 177578 400294 177648 400350
rect 177328 400226 177648 400294
rect 177328 400170 177398 400226
rect 177454 400170 177522 400226
rect 177578 400170 177648 400226
rect 177328 400102 177648 400170
rect 177328 400046 177398 400102
rect 177454 400046 177522 400102
rect 177578 400046 177648 400102
rect 177328 399978 177648 400046
rect 177328 399922 177398 399978
rect 177454 399922 177522 399978
rect 177578 399922 177648 399978
rect 177328 399888 177648 399922
rect 208048 400350 208368 400384
rect 208048 400294 208118 400350
rect 208174 400294 208242 400350
rect 208298 400294 208368 400350
rect 208048 400226 208368 400294
rect 208048 400170 208118 400226
rect 208174 400170 208242 400226
rect 208298 400170 208368 400226
rect 208048 400102 208368 400170
rect 208048 400046 208118 400102
rect 208174 400046 208242 400102
rect 208298 400046 208368 400102
rect 208048 399978 208368 400046
rect 208048 399922 208118 399978
rect 208174 399922 208242 399978
rect 208298 399922 208368 399978
rect 208048 399888 208368 399922
rect 238768 400350 239088 400384
rect 238768 400294 238838 400350
rect 238894 400294 238962 400350
rect 239018 400294 239088 400350
rect 238768 400226 239088 400294
rect 238768 400170 238838 400226
rect 238894 400170 238962 400226
rect 239018 400170 239088 400226
rect 238768 400102 239088 400170
rect 238768 400046 238838 400102
rect 238894 400046 238962 400102
rect 239018 400046 239088 400102
rect 238768 399978 239088 400046
rect 238768 399922 238838 399978
rect 238894 399922 238962 399978
rect 239018 399922 239088 399978
rect 238768 399888 239088 399922
rect 269488 400350 269808 400384
rect 269488 400294 269558 400350
rect 269614 400294 269682 400350
rect 269738 400294 269808 400350
rect 269488 400226 269808 400294
rect 269488 400170 269558 400226
rect 269614 400170 269682 400226
rect 269738 400170 269808 400226
rect 269488 400102 269808 400170
rect 269488 400046 269558 400102
rect 269614 400046 269682 400102
rect 269738 400046 269808 400102
rect 269488 399978 269808 400046
rect 269488 399922 269558 399978
rect 269614 399922 269682 399978
rect 269738 399922 269808 399978
rect 269488 399888 269808 399922
rect 300208 400350 300528 400384
rect 300208 400294 300278 400350
rect 300334 400294 300402 400350
rect 300458 400294 300528 400350
rect 300208 400226 300528 400294
rect 300208 400170 300278 400226
rect 300334 400170 300402 400226
rect 300458 400170 300528 400226
rect 300208 400102 300528 400170
rect 300208 400046 300278 400102
rect 300334 400046 300402 400102
rect 300458 400046 300528 400102
rect 300208 399978 300528 400046
rect 300208 399922 300278 399978
rect 300334 399922 300402 399978
rect 300458 399922 300528 399978
rect 300208 399888 300528 399922
rect 330928 400350 331248 400384
rect 330928 400294 330998 400350
rect 331054 400294 331122 400350
rect 331178 400294 331248 400350
rect 330928 400226 331248 400294
rect 330928 400170 330998 400226
rect 331054 400170 331122 400226
rect 331178 400170 331248 400226
rect 330928 400102 331248 400170
rect 330928 400046 330998 400102
rect 331054 400046 331122 400102
rect 331178 400046 331248 400102
rect 330928 399978 331248 400046
rect 330928 399922 330998 399978
rect 331054 399922 331122 399978
rect 331178 399922 331248 399978
rect 330928 399888 331248 399922
rect 361648 400350 361968 400384
rect 361648 400294 361718 400350
rect 361774 400294 361842 400350
rect 361898 400294 361968 400350
rect 361648 400226 361968 400294
rect 361648 400170 361718 400226
rect 361774 400170 361842 400226
rect 361898 400170 361968 400226
rect 361648 400102 361968 400170
rect 361648 400046 361718 400102
rect 361774 400046 361842 400102
rect 361898 400046 361968 400102
rect 361648 399978 361968 400046
rect 361648 399922 361718 399978
rect 361774 399922 361842 399978
rect 361898 399922 361968 399978
rect 361648 399888 361968 399922
rect 392368 400350 392688 400384
rect 392368 400294 392438 400350
rect 392494 400294 392562 400350
rect 392618 400294 392688 400350
rect 392368 400226 392688 400294
rect 392368 400170 392438 400226
rect 392494 400170 392562 400226
rect 392618 400170 392688 400226
rect 392368 400102 392688 400170
rect 392368 400046 392438 400102
rect 392494 400046 392562 400102
rect 392618 400046 392688 400102
rect 392368 399978 392688 400046
rect 392368 399922 392438 399978
rect 392494 399922 392562 399978
rect 392618 399922 392688 399978
rect 392368 399888 392688 399922
rect 423088 400350 423408 400384
rect 423088 400294 423158 400350
rect 423214 400294 423282 400350
rect 423338 400294 423408 400350
rect 423088 400226 423408 400294
rect 423088 400170 423158 400226
rect 423214 400170 423282 400226
rect 423338 400170 423408 400226
rect 423088 400102 423408 400170
rect 423088 400046 423158 400102
rect 423214 400046 423282 400102
rect 423338 400046 423408 400102
rect 423088 399978 423408 400046
rect 423088 399922 423158 399978
rect 423214 399922 423282 399978
rect 423338 399922 423408 399978
rect 423088 399888 423408 399922
rect 453808 400350 454128 400384
rect 453808 400294 453878 400350
rect 453934 400294 454002 400350
rect 454058 400294 454128 400350
rect 453808 400226 454128 400294
rect 453808 400170 453878 400226
rect 453934 400170 454002 400226
rect 454058 400170 454128 400226
rect 453808 400102 454128 400170
rect 453808 400046 453878 400102
rect 453934 400046 454002 400102
rect 454058 400046 454128 400102
rect 453808 399978 454128 400046
rect 453808 399922 453878 399978
rect 453934 399922 454002 399978
rect 454058 399922 454128 399978
rect 453808 399888 454128 399922
rect 484528 400350 484848 400384
rect 484528 400294 484598 400350
rect 484654 400294 484722 400350
rect 484778 400294 484848 400350
rect 484528 400226 484848 400294
rect 484528 400170 484598 400226
rect 484654 400170 484722 400226
rect 484778 400170 484848 400226
rect 484528 400102 484848 400170
rect 484528 400046 484598 400102
rect 484654 400046 484722 400102
rect 484778 400046 484848 400102
rect 484528 399978 484848 400046
rect 484528 399922 484598 399978
rect 484654 399922 484722 399978
rect 484778 399922 484848 399978
rect 484528 399888 484848 399922
rect 515248 400350 515568 400384
rect 515248 400294 515318 400350
rect 515374 400294 515442 400350
rect 515498 400294 515568 400350
rect 515248 400226 515568 400294
rect 515248 400170 515318 400226
rect 515374 400170 515442 400226
rect 515498 400170 515568 400226
rect 515248 400102 515568 400170
rect 515248 400046 515318 400102
rect 515374 400046 515442 400102
rect 515498 400046 515568 400102
rect 515248 399978 515568 400046
rect 515248 399922 515318 399978
rect 515374 399922 515442 399978
rect 515498 399922 515568 399978
rect 515248 399888 515568 399922
rect 545968 400350 546288 400384
rect 545968 400294 546038 400350
rect 546094 400294 546162 400350
rect 546218 400294 546288 400350
rect 545968 400226 546288 400294
rect 545968 400170 546038 400226
rect 546094 400170 546162 400226
rect 546218 400170 546288 400226
rect 545968 400102 546288 400170
rect 545968 400046 546038 400102
rect 546094 400046 546162 400102
rect 546218 400046 546288 400102
rect 545968 399978 546288 400046
rect 545968 399922 546038 399978
rect 546094 399922 546162 399978
rect 546218 399922 546288 399978
rect 545968 399888 546288 399922
rect 561154 400350 561774 417922
rect 561154 400294 561250 400350
rect 561306 400294 561374 400350
rect 561430 400294 561498 400350
rect 561554 400294 561622 400350
rect 561678 400294 561774 400350
rect 561154 400226 561774 400294
rect 561154 400170 561250 400226
rect 561306 400170 561374 400226
rect 561430 400170 561498 400226
rect 561554 400170 561622 400226
rect 561678 400170 561774 400226
rect 561154 400102 561774 400170
rect 561154 400046 561250 400102
rect 561306 400046 561374 400102
rect 561430 400046 561498 400102
rect 561554 400046 561622 400102
rect 561678 400046 561774 400102
rect 561154 399978 561774 400046
rect 561154 399922 561250 399978
rect 561306 399922 561374 399978
rect 561430 399922 561498 399978
rect 561554 399922 561622 399978
rect 561678 399922 561774 399978
rect 131248 388350 131568 388384
rect 131248 388294 131318 388350
rect 131374 388294 131442 388350
rect 131498 388294 131568 388350
rect 131248 388226 131568 388294
rect 131248 388170 131318 388226
rect 131374 388170 131442 388226
rect 131498 388170 131568 388226
rect 131248 388102 131568 388170
rect 131248 388046 131318 388102
rect 131374 388046 131442 388102
rect 131498 388046 131568 388102
rect 131248 387978 131568 388046
rect 131248 387922 131318 387978
rect 131374 387922 131442 387978
rect 131498 387922 131568 387978
rect 131248 387888 131568 387922
rect 161968 388350 162288 388384
rect 161968 388294 162038 388350
rect 162094 388294 162162 388350
rect 162218 388294 162288 388350
rect 161968 388226 162288 388294
rect 161968 388170 162038 388226
rect 162094 388170 162162 388226
rect 162218 388170 162288 388226
rect 161968 388102 162288 388170
rect 161968 388046 162038 388102
rect 162094 388046 162162 388102
rect 162218 388046 162288 388102
rect 161968 387978 162288 388046
rect 161968 387922 162038 387978
rect 162094 387922 162162 387978
rect 162218 387922 162288 387978
rect 161968 387888 162288 387922
rect 192688 388350 193008 388384
rect 192688 388294 192758 388350
rect 192814 388294 192882 388350
rect 192938 388294 193008 388350
rect 192688 388226 193008 388294
rect 192688 388170 192758 388226
rect 192814 388170 192882 388226
rect 192938 388170 193008 388226
rect 192688 388102 193008 388170
rect 192688 388046 192758 388102
rect 192814 388046 192882 388102
rect 192938 388046 193008 388102
rect 192688 387978 193008 388046
rect 192688 387922 192758 387978
rect 192814 387922 192882 387978
rect 192938 387922 193008 387978
rect 192688 387888 193008 387922
rect 223408 388350 223728 388384
rect 223408 388294 223478 388350
rect 223534 388294 223602 388350
rect 223658 388294 223728 388350
rect 223408 388226 223728 388294
rect 223408 388170 223478 388226
rect 223534 388170 223602 388226
rect 223658 388170 223728 388226
rect 223408 388102 223728 388170
rect 223408 388046 223478 388102
rect 223534 388046 223602 388102
rect 223658 388046 223728 388102
rect 223408 387978 223728 388046
rect 223408 387922 223478 387978
rect 223534 387922 223602 387978
rect 223658 387922 223728 387978
rect 223408 387888 223728 387922
rect 254128 388350 254448 388384
rect 254128 388294 254198 388350
rect 254254 388294 254322 388350
rect 254378 388294 254448 388350
rect 254128 388226 254448 388294
rect 254128 388170 254198 388226
rect 254254 388170 254322 388226
rect 254378 388170 254448 388226
rect 254128 388102 254448 388170
rect 254128 388046 254198 388102
rect 254254 388046 254322 388102
rect 254378 388046 254448 388102
rect 254128 387978 254448 388046
rect 254128 387922 254198 387978
rect 254254 387922 254322 387978
rect 254378 387922 254448 387978
rect 254128 387888 254448 387922
rect 284848 388350 285168 388384
rect 284848 388294 284918 388350
rect 284974 388294 285042 388350
rect 285098 388294 285168 388350
rect 284848 388226 285168 388294
rect 284848 388170 284918 388226
rect 284974 388170 285042 388226
rect 285098 388170 285168 388226
rect 284848 388102 285168 388170
rect 284848 388046 284918 388102
rect 284974 388046 285042 388102
rect 285098 388046 285168 388102
rect 284848 387978 285168 388046
rect 284848 387922 284918 387978
rect 284974 387922 285042 387978
rect 285098 387922 285168 387978
rect 284848 387888 285168 387922
rect 315568 388350 315888 388384
rect 315568 388294 315638 388350
rect 315694 388294 315762 388350
rect 315818 388294 315888 388350
rect 315568 388226 315888 388294
rect 315568 388170 315638 388226
rect 315694 388170 315762 388226
rect 315818 388170 315888 388226
rect 315568 388102 315888 388170
rect 315568 388046 315638 388102
rect 315694 388046 315762 388102
rect 315818 388046 315888 388102
rect 315568 387978 315888 388046
rect 315568 387922 315638 387978
rect 315694 387922 315762 387978
rect 315818 387922 315888 387978
rect 315568 387888 315888 387922
rect 346288 388350 346608 388384
rect 346288 388294 346358 388350
rect 346414 388294 346482 388350
rect 346538 388294 346608 388350
rect 346288 388226 346608 388294
rect 346288 388170 346358 388226
rect 346414 388170 346482 388226
rect 346538 388170 346608 388226
rect 346288 388102 346608 388170
rect 346288 388046 346358 388102
rect 346414 388046 346482 388102
rect 346538 388046 346608 388102
rect 346288 387978 346608 388046
rect 346288 387922 346358 387978
rect 346414 387922 346482 387978
rect 346538 387922 346608 387978
rect 346288 387888 346608 387922
rect 377008 388350 377328 388384
rect 377008 388294 377078 388350
rect 377134 388294 377202 388350
rect 377258 388294 377328 388350
rect 377008 388226 377328 388294
rect 377008 388170 377078 388226
rect 377134 388170 377202 388226
rect 377258 388170 377328 388226
rect 377008 388102 377328 388170
rect 377008 388046 377078 388102
rect 377134 388046 377202 388102
rect 377258 388046 377328 388102
rect 377008 387978 377328 388046
rect 377008 387922 377078 387978
rect 377134 387922 377202 387978
rect 377258 387922 377328 387978
rect 377008 387888 377328 387922
rect 407728 388350 408048 388384
rect 407728 388294 407798 388350
rect 407854 388294 407922 388350
rect 407978 388294 408048 388350
rect 407728 388226 408048 388294
rect 407728 388170 407798 388226
rect 407854 388170 407922 388226
rect 407978 388170 408048 388226
rect 407728 388102 408048 388170
rect 407728 388046 407798 388102
rect 407854 388046 407922 388102
rect 407978 388046 408048 388102
rect 407728 387978 408048 388046
rect 407728 387922 407798 387978
rect 407854 387922 407922 387978
rect 407978 387922 408048 387978
rect 407728 387888 408048 387922
rect 438448 388350 438768 388384
rect 438448 388294 438518 388350
rect 438574 388294 438642 388350
rect 438698 388294 438768 388350
rect 438448 388226 438768 388294
rect 438448 388170 438518 388226
rect 438574 388170 438642 388226
rect 438698 388170 438768 388226
rect 438448 388102 438768 388170
rect 438448 388046 438518 388102
rect 438574 388046 438642 388102
rect 438698 388046 438768 388102
rect 438448 387978 438768 388046
rect 438448 387922 438518 387978
rect 438574 387922 438642 387978
rect 438698 387922 438768 387978
rect 438448 387888 438768 387922
rect 469168 388350 469488 388384
rect 469168 388294 469238 388350
rect 469294 388294 469362 388350
rect 469418 388294 469488 388350
rect 469168 388226 469488 388294
rect 469168 388170 469238 388226
rect 469294 388170 469362 388226
rect 469418 388170 469488 388226
rect 469168 388102 469488 388170
rect 469168 388046 469238 388102
rect 469294 388046 469362 388102
rect 469418 388046 469488 388102
rect 469168 387978 469488 388046
rect 469168 387922 469238 387978
rect 469294 387922 469362 387978
rect 469418 387922 469488 387978
rect 469168 387888 469488 387922
rect 499888 388350 500208 388384
rect 499888 388294 499958 388350
rect 500014 388294 500082 388350
rect 500138 388294 500208 388350
rect 499888 388226 500208 388294
rect 499888 388170 499958 388226
rect 500014 388170 500082 388226
rect 500138 388170 500208 388226
rect 499888 388102 500208 388170
rect 499888 388046 499958 388102
rect 500014 388046 500082 388102
rect 500138 388046 500208 388102
rect 499888 387978 500208 388046
rect 499888 387922 499958 387978
rect 500014 387922 500082 387978
rect 500138 387922 500208 387978
rect 499888 387888 500208 387922
rect 530608 388350 530928 388384
rect 530608 388294 530678 388350
rect 530734 388294 530802 388350
rect 530858 388294 530928 388350
rect 530608 388226 530928 388294
rect 530608 388170 530678 388226
rect 530734 388170 530802 388226
rect 530858 388170 530928 388226
rect 530608 388102 530928 388170
rect 530608 388046 530678 388102
rect 530734 388046 530802 388102
rect 530858 388046 530928 388102
rect 530608 387978 530928 388046
rect 530608 387922 530678 387978
rect 530734 387922 530802 387978
rect 530858 387922 530928 387978
rect 530608 387888 530928 387922
rect 111154 382294 111250 382350
rect 111306 382294 111374 382350
rect 111430 382294 111498 382350
rect 111554 382294 111622 382350
rect 111678 382294 111774 382350
rect 111154 382226 111774 382294
rect 111154 382170 111250 382226
rect 111306 382170 111374 382226
rect 111430 382170 111498 382226
rect 111554 382170 111622 382226
rect 111678 382170 111774 382226
rect 111154 382102 111774 382170
rect 111154 382046 111250 382102
rect 111306 382046 111374 382102
rect 111430 382046 111498 382102
rect 111554 382046 111622 382102
rect 111678 382046 111774 382102
rect 111154 381978 111774 382046
rect 111154 381922 111250 381978
rect 111306 381922 111374 381978
rect 111430 381922 111498 381978
rect 111554 381922 111622 381978
rect 111678 381922 111774 381978
rect 96874 370294 96970 370350
rect 97026 370294 97094 370350
rect 97150 370294 97218 370350
rect 97274 370294 97342 370350
rect 97398 370294 97494 370350
rect 96874 370226 97494 370294
rect 96874 370170 96970 370226
rect 97026 370170 97094 370226
rect 97150 370170 97218 370226
rect 97274 370170 97342 370226
rect 97398 370170 97494 370226
rect 96874 370102 97494 370170
rect 96874 370046 96970 370102
rect 97026 370046 97094 370102
rect 97150 370046 97218 370102
rect 97274 370046 97342 370102
rect 97398 370046 97494 370102
rect 96874 369978 97494 370046
rect 96874 369922 96970 369978
rect 97026 369922 97094 369978
rect 97150 369922 97218 369978
rect 97274 369922 97342 369978
rect 97398 369922 97494 369978
rect 96874 352350 97494 369922
rect 100528 370350 100848 370384
rect 100528 370294 100598 370350
rect 100654 370294 100722 370350
rect 100778 370294 100848 370350
rect 100528 370226 100848 370294
rect 100528 370170 100598 370226
rect 100654 370170 100722 370226
rect 100778 370170 100848 370226
rect 100528 370102 100848 370170
rect 100528 370046 100598 370102
rect 100654 370046 100722 370102
rect 100778 370046 100848 370102
rect 100528 369978 100848 370046
rect 100528 369922 100598 369978
rect 100654 369922 100722 369978
rect 100778 369922 100848 369978
rect 100528 369888 100848 369922
rect 111154 364350 111774 381922
rect 115888 382350 116208 382384
rect 115888 382294 115958 382350
rect 116014 382294 116082 382350
rect 116138 382294 116208 382350
rect 115888 382226 116208 382294
rect 115888 382170 115958 382226
rect 116014 382170 116082 382226
rect 116138 382170 116208 382226
rect 115888 382102 116208 382170
rect 115888 382046 115958 382102
rect 116014 382046 116082 382102
rect 116138 382046 116208 382102
rect 115888 381978 116208 382046
rect 115888 381922 115958 381978
rect 116014 381922 116082 381978
rect 116138 381922 116208 381978
rect 115888 381888 116208 381922
rect 146608 382350 146928 382384
rect 146608 382294 146678 382350
rect 146734 382294 146802 382350
rect 146858 382294 146928 382350
rect 146608 382226 146928 382294
rect 146608 382170 146678 382226
rect 146734 382170 146802 382226
rect 146858 382170 146928 382226
rect 146608 382102 146928 382170
rect 146608 382046 146678 382102
rect 146734 382046 146802 382102
rect 146858 382046 146928 382102
rect 146608 381978 146928 382046
rect 146608 381922 146678 381978
rect 146734 381922 146802 381978
rect 146858 381922 146928 381978
rect 146608 381888 146928 381922
rect 177328 382350 177648 382384
rect 177328 382294 177398 382350
rect 177454 382294 177522 382350
rect 177578 382294 177648 382350
rect 177328 382226 177648 382294
rect 177328 382170 177398 382226
rect 177454 382170 177522 382226
rect 177578 382170 177648 382226
rect 177328 382102 177648 382170
rect 177328 382046 177398 382102
rect 177454 382046 177522 382102
rect 177578 382046 177648 382102
rect 177328 381978 177648 382046
rect 177328 381922 177398 381978
rect 177454 381922 177522 381978
rect 177578 381922 177648 381978
rect 177328 381888 177648 381922
rect 208048 382350 208368 382384
rect 208048 382294 208118 382350
rect 208174 382294 208242 382350
rect 208298 382294 208368 382350
rect 208048 382226 208368 382294
rect 208048 382170 208118 382226
rect 208174 382170 208242 382226
rect 208298 382170 208368 382226
rect 208048 382102 208368 382170
rect 208048 382046 208118 382102
rect 208174 382046 208242 382102
rect 208298 382046 208368 382102
rect 208048 381978 208368 382046
rect 208048 381922 208118 381978
rect 208174 381922 208242 381978
rect 208298 381922 208368 381978
rect 208048 381888 208368 381922
rect 238768 382350 239088 382384
rect 238768 382294 238838 382350
rect 238894 382294 238962 382350
rect 239018 382294 239088 382350
rect 238768 382226 239088 382294
rect 238768 382170 238838 382226
rect 238894 382170 238962 382226
rect 239018 382170 239088 382226
rect 238768 382102 239088 382170
rect 238768 382046 238838 382102
rect 238894 382046 238962 382102
rect 239018 382046 239088 382102
rect 238768 381978 239088 382046
rect 238768 381922 238838 381978
rect 238894 381922 238962 381978
rect 239018 381922 239088 381978
rect 238768 381888 239088 381922
rect 269488 382350 269808 382384
rect 269488 382294 269558 382350
rect 269614 382294 269682 382350
rect 269738 382294 269808 382350
rect 269488 382226 269808 382294
rect 269488 382170 269558 382226
rect 269614 382170 269682 382226
rect 269738 382170 269808 382226
rect 269488 382102 269808 382170
rect 269488 382046 269558 382102
rect 269614 382046 269682 382102
rect 269738 382046 269808 382102
rect 269488 381978 269808 382046
rect 269488 381922 269558 381978
rect 269614 381922 269682 381978
rect 269738 381922 269808 381978
rect 269488 381888 269808 381922
rect 300208 382350 300528 382384
rect 300208 382294 300278 382350
rect 300334 382294 300402 382350
rect 300458 382294 300528 382350
rect 300208 382226 300528 382294
rect 300208 382170 300278 382226
rect 300334 382170 300402 382226
rect 300458 382170 300528 382226
rect 300208 382102 300528 382170
rect 300208 382046 300278 382102
rect 300334 382046 300402 382102
rect 300458 382046 300528 382102
rect 300208 381978 300528 382046
rect 300208 381922 300278 381978
rect 300334 381922 300402 381978
rect 300458 381922 300528 381978
rect 300208 381888 300528 381922
rect 330928 382350 331248 382384
rect 330928 382294 330998 382350
rect 331054 382294 331122 382350
rect 331178 382294 331248 382350
rect 330928 382226 331248 382294
rect 330928 382170 330998 382226
rect 331054 382170 331122 382226
rect 331178 382170 331248 382226
rect 330928 382102 331248 382170
rect 330928 382046 330998 382102
rect 331054 382046 331122 382102
rect 331178 382046 331248 382102
rect 330928 381978 331248 382046
rect 330928 381922 330998 381978
rect 331054 381922 331122 381978
rect 331178 381922 331248 381978
rect 330928 381888 331248 381922
rect 361648 382350 361968 382384
rect 361648 382294 361718 382350
rect 361774 382294 361842 382350
rect 361898 382294 361968 382350
rect 361648 382226 361968 382294
rect 361648 382170 361718 382226
rect 361774 382170 361842 382226
rect 361898 382170 361968 382226
rect 361648 382102 361968 382170
rect 361648 382046 361718 382102
rect 361774 382046 361842 382102
rect 361898 382046 361968 382102
rect 361648 381978 361968 382046
rect 361648 381922 361718 381978
rect 361774 381922 361842 381978
rect 361898 381922 361968 381978
rect 361648 381888 361968 381922
rect 392368 382350 392688 382384
rect 392368 382294 392438 382350
rect 392494 382294 392562 382350
rect 392618 382294 392688 382350
rect 392368 382226 392688 382294
rect 392368 382170 392438 382226
rect 392494 382170 392562 382226
rect 392618 382170 392688 382226
rect 392368 382102 392688 382170
rect 392368 382046 392438 382102
rect 392494 382046 392562 382102
rect 392618 382046 392688 382102
rect 392368 381978 392688 382046
rect 392368 381922 392438 381978
rect 392494 381922 392562 381978
rect 392618 381922 392688 381978
rect 392368 381888 392688 381922
rect 423088 382350 423408 382384
rect 423088 382294 423158 382350
rect 423214 382294 423282 382350
rect 423338 382294 423408 382350
rect 423088 382226 423408 382294
rect 423088 382170 423158 382226
rect 423214 382170 423282 382226
rect 423338 382170 423408 382226
rect 423088 382102 423408 382170
rect 423088 382046 423158 382102
rect 423214 382046 423282 382102
rect 423338 382046 423408 382102
rect 423088 381978 423408 382046
rect 423088 381922 423158 381978
rect 423214 381922 423282 381978
rect 423338 381922 423408 381978
rect 423088 381888 423408 381922
rect 453808 382350 454128 382384
rect 453808 382294 453878 382350
rect 453934 382294 454002 382350
rect 454058 382294 454128 382350
rect 453808 382226 454128 382294
rect 453808 382170 453878 382226
rect 453934 382170 454002 382226
rect 454058 382170 454128 382226
rect 453808 382102 454128 382170
rect 453808 382046 453878 382102
rect 453934 382046 454002 382102
rect 454058 382046 454128 382102
rect 453808 381978 454128 382046
rect 453808 381922 453878 381978
rect 453934 381922 454002 381978
rect 454058 381922 454128 381978
rect 453808 381888 454128 381922
rect 484528 382350 484848 382384
rect 484528 382294 484598 382350
rect 484654 382294 484722 382350
rect 484778 382294 484848 382350
rect 484528 382226 484848 382294
rect 484528 382170 484598 382226
rect 484654 382170 484722 382226
rect 484778 382170 484848 382226
rect 484528 382102 484848 382170
rect 484528 382046 484598 382102
rect 484654 382046 484722 382102
rect 484778 382046 484848 382102
rect 484528 381978 484848 382046
rect 484528 381922 484598 381978
rect 484654 381922 484722 381978
rect 484778 381922 484848 381978
rect 484528 381888 484848 381922
rect 515248 382350 515568 382384
rect 515248 382294 515318 382350
rect 515374 382294 515442 382350
rect 515498 382294 515568 382350
rect 515248 382226 515568 382294
rect 515248 382170 515318 382226
rect 515374 382170 515442 382226
rect 515498 382170 515568 382226
rect 515248 382102 515568 382170
rect 515248 382046 515318 382102
rect 515374 382046 515442 382102
rect 515498 382046 515568 382102
rect 515248 381978 515568 382046
rect 515248 381922 515318 381978
rect 515374 381922 515442 381978
rect 515498 381922 515568 381978
rect 515248 381888 515568 381922
rect 545968 382350 546288 382384
rect 545968 382294 546038 382350
rect 546094 382294 546162 382350
rect 546218 382294 546288 382350
rect 545968 382226 546288 382294
rect 545968 382170 546038 382226
rect 546094 382170 546162 382226
rect 546218 382170 546288 382226
rect 545968 382102 546288 382170
rect 545968 382046 546038 382102
rect 546094 382046 546162 382102
rect 546218 382046 546288 382102
rect 545968 381978 546288 382046
rect 545968 381922 546038 381978
rect 546094 381922 546162 381978
rect 546218 381922 546288 381978
rect 545968 381888 546288 381922
rect 561154 382350 561774 399922
rect 561154 382294 561250 382350
rect 561306 382294 561374 382350
rect 561430 382294 561498 382350
rect 561554 382294 561622 382350
rect 561678 382294 561774 382350
rect 561154 382226 561774 382294
rect 561154 382170 561250 382226
rect 561306 382170 561374 382226
rect 561430 382170 561498 382226
rect 561554 382170 561622 382226
rect 561678 382170 561774 382226
rect 561154 382102 561774 382170
rect 561154 382046 561250 382102
rect 561306 382046 561374 382102
rect 561430 382046 561498 382102
rect 561554 382046 561622 382102
rect 561678 382046 561774 382102
rect 561154 381978 561774 382046
rect 561154 381922 561250 381978
rect 561306 381922 561374 381978
rect 561430 381922 561498 381978
rect 561554 381922 561622 381978
rect 561678 381922 561774 381978
rect 131248 370350 131568 370384
rect 131248 370294 131318 370350
rect 131374 370294 131442 370350
rect 131498 370294 131568 370350
rect 131248 370226 131568 370294
rect 131248 370170 131318 370226
rect 131374 370170 131442 370226
rect 131498 370170 131568 370226
rect 131248 370102 131568 370170
rect 131248 370046 131318 370102
rect 131374 370046 131442 370102
rect 131498 370046 131568 370102
rect 131248 369978 131568 370046
rect 131248 369922 131318 369978
rect 131374 369922 131442 369978
rect 131498 369922 131568 369978
rect 131248 369888 131568 369922
rect 161968 370350 162288 370384
rect 161968 370294 162038 370350
rect 162094 370294 162162 370350
rect 162218 370294 162288 370350
rect 161968 370226 162288 370294
rect 161968 370170 162038 370226
rect 162094 370170 162162 370226
rect 162218 370170 162288 370226
rect 161968 370102 162288 370170
rect 161968 370046 162038 370102
rect 162094 370046 162162 370102
rect 162218 370046 162288 370102
rect 161968 369978 162288 370046
rect 161968 369922 162038 369978
rect 162094 369922 162162 369978
rect 162218 369922 162288 369978
rect 161968 369888 162288 369922
rect 192688 370350 193008 370384
rect 192688 370294 192758 370350
rect 192814 370294 192882 370350
rect 192938 370294 193008 370350
rect 192688 370226 193008 370294
rect 192688 370170 192758 370226
rect 192814 370170 192882 370226
rect 192938 370170 193008 370226
rect 192688 370102 193008 370170
rect 192688 370046 192758 370102
rect 192814 370046 192882 370102
rect 192938 370046 193008 370102
rect 192688 369978 193008 370046
rect 192688 369922 192758 369978
rect 192814 369922 192882 369978
rect 192938 369922 193008 369978
rect 192688 369888 193008 369922
rect 223408 370350 223728 370384
rect 223408 370294 223478 370350
rect 223534 370294 223602 370350
rect 223658 370294 223728 370350
rect 223408 370226 223728 370294
rect 223408 370170 223478 370226
rect 223534 370170 223602 370226
rect 223658 370170 223728 370226
rect 223408 370102 223728 370170
rect 223408 370046 223478 370102
rect 223534 370046 223602 370102
rect 223658 370046 223728 370102
rect 223408 369978 223728 370046
rect 223408 369922 223478 369978
rect 223534 369922 223602 369978
rect 223658 369922 223728 369978
rect 223408 369888 223728 369922
rect 254128 370350 254448 370384
rect 254128 370294 254198 370350
rect 254254 370294 254322 370350
rect 254378 370294 254448 370350
rect 254128 370226 254448 370294
rect 254128 370170 254198 370226
rect 254254 370170 254322 370226
rect 254378 370170 254448 370226
rect 254128 370102 254448 370170
rect 254128 370046 254198 370102
rect 254254 370046 254322 370102
rect 254378 370046 254448 370102
rect 254128 369978 254448 370046
rect 254128 369922 254198 369978
rect 254254 369922 254322 369978
rect 254378 369922 254448 369978
rect 254128 369888 254448 369922
rect 284848 370350 285168 370384
rect 284848 370294 284918 370350
rect 284974 370294 285042 370350
rect 285098 370294 285168 370350
rect 284848 370226 285168 370294
rect 284848 370170 284918 370226
rect 284974 370170 285042 370226
rect 285098 370170 285168 370226
rect 284848 370102 285168 370170
rect 284848 370046 284918 370102
rect 284974 370046 285042 370102
rect 285098 370046 285168 370102
rect 284848 369978 285168 370046
rect 284848 369922 284918 369978
rect 284974 369922 285042 369978
rect 285098 369922 285168 369978
rect 284848 369888 285168 369922
rect 315568 370350 315888 370384
rect 315568 370294 315638 370350
rect 315694 370294 315762 370350
rect 315818 370294 315888 370350
rect 315568 370226 315888 370294
rect 315568 370170 315638 370226
rect 315694 370170 315762 370226
rect 315818 370170 315888 370226
rect 315568 370102 315888 370170
rect 315568 370046 315638 370102
rect 315694 370046 315762 370102
rect 315818 370046 315888 370102
rect 315568 369978 315888 370046
rect 315568 369922 315638 369978
rect 315694 369922 315762 369978
rect 315818 369922 315888 369978
rect 315568 369888 315888 369922
rect 346288 370350 346608 370384
rect 346288 370294 346358 370350
rect 346414 370294 346482 370350
rect 346538 370294 346608 370350
rect 346288 370226 346608 370294
rect 346288 370170 346358 370226
rect 346414 370170 346482 370226
rect 346538 370170 346608 370226
rect 346288 370102 346608 370170
rect 346288 370046 346358 370102
rect 346414 370046 346482 370102
rect 346538 370046 346608 370102
rect 346288 369978 346608 370046
rect 346288 369922 346358 369978
rect 346414 369922 346482 369978
rect 346538 369922 346608 369978
rect 346288 369888 346608 369922
rect 377008 370350 377328 370384
rect 377008 370294 377078 370350
rect 377134 370294 377202 370350
rect 377258 370294 377328 370350
rect 377008 370226 377328 370294
rect 377008 370170 377078 370226
rect 377134 370170 377202 370226
rect 377258 370170 377328 370226
rect 377008 370102 377328 370170
rect 377008 370046 377078 370102
rect 377134 370046 377202 370102
rect 377258 370046 377328 370102
rect 377008 369978 377328 370046
rect 377008 369922 377078 369978
rect 377134 369922 377202 369978
rect 377258 369922 377328 369978
rect 377008 369888 377328 369922
rect 407728 370350 408048 370384
rect 407728 370294 407798 370350
rect 407854 370294 407922 370350
rect 407978 370294 408048 370350
rect 407728 370226 408048 370294
rect 407728 370170 407798 370226
rect 407854 370170 407922 370226
rect 407978 370170 408048 370226
rect 407728 370102 408048 370170
rect 407728 370046 407798 370102
rect 407854 370046 407922 370102
rect 407978 370046 408048 370102
rect 407728 369978 408048 370046
rect 407728 369922 407798 369978
rect 407854 369922 407922 369978
rect 407978 369922 408048 369978
rect 407728 369888 408048 369922
rect 438448 370350 438768 370384
rect 438448 370294 438518 370350
rect 438574 370294 438642 370350
rect 438698 370294 438768 370350
rect 438448 370226 438768 370294
rect 438448 370170 438518 370226
rect 438574 370170 438642 370226
rect 438698 370170 438768 370226
rect 438448 370102 438768 370170
rect 438448 370046 438518 370102
rect 438574 370046 438642 370102
rect 438698 370046 438768 370102
rect 438448 369978 438768 370046
rect 438448 369922 438518 369978
rect 438574 369922 438642 369978
rect 438698 369922 438768 369978
rect 438448 369888 438768 369922
rect 469168 370350 469488 370384
rect 469168 370294 469238 370350
rect 469294 370294 469362 370350
rect 469418 370294 469488 370350
rect 469168 370226 469488 370294
rect 469168 370170 469238 370226
rect 469294 370170 469362 370226
rect 469418 370170 469488 370226
rect 469168 370102 469488 370170
rect 469168 370046 469238 370102
rect 469294 370046 469362 370102
rect 469418 370046 469488 370102
rect 469168 369978 469488 370046
rect 469168 369922 469238 369978
rect 469294 369922 469362 369978
rect 469418 369922 469488 369978
rect 469168 369888 469488 369922
rect 499888 370350 500208 370384
rect 499888 370294 499958 370350
rect 500014 370294 500082 370350
rect 500138 370294 500208 370350
rect 499888 370226 500208 370294
rect 499888 370170 499958 370226
rect 500014 370170 500082 370226
rect 500138 370170 500208 370226
rect 499888 370102 500208 370170
rect 499888 370046 499958 370102
rect 500014 370046 500082 370102
rect 500138 370046 500208 370102
rect 499888 369978 500208 370046
rect 499888 369922 499958 369978
rect 500014 369922 500082 369978
rect 500138 369922 500208 369978
rect 499888 369888 500208 369922
rect 530608 370350 530928 370384
rect 530608 370294 530678 370350
rect 530734 370294 530802 370350
rect 530858 370294 530928 370350
rect 530608 370226 530928 370294
rect 530608 370170 530678 370226
rect 530734 370170 530802 370226
rect 530858 370170 530928 370226
rect 530608 370102 530928 370170
rect 530608 370046 530678 370102
rect 530734 370046 530802 370102
rect 530858 370046 530928 370102
rect 530608 369978 530928 370046
rect 530608 369922 530678 369978
rect 530734 369922 530802 369978
rect 530858 369922 530928 369978
rect 530608 369888 530928 369922
rect 111154 364294 111250 364350
rect 111306 364294 111374 364350
rect 111430 364294 111498 364350
rect 111554 364294 111622 364350
rect 111678 364294 111774 364350
rect 111154 364226 111774 364294
rect 111154 364170 111250 364226
rect 111306 364170 111374 364226
rect 111430 364170 111498 364226
rect 111554 364170 111622 364226
rect 111678 364170 111774 364226
rect 111154 364102 111774 364170
rect 111154 364046 111250 364102
rect 111306 364046 111374 364102
rect 111430 364046 111498 364102
rect 111554 364046 111622 364102
rect 111678 364046 111774 364102
rect 111154 363978 111774 364046
rect 111154 363922 111250 363978
rect 111306 363922 111374 363978
rect 111430 363922 111498 363978
rect 111554 363922 111622 363978
rect 111678 363922 111774 363978
rect 96874 352294 96970 352350
rect 97026 352294 97094 352350
rect 97150 352294 97218 352350
rect 97274 352294 97342 352350
rect 97398 352294 97494 352350
rect 96874 352226 97494 352294
rect 96874 352170 96970 352226
rect 97026 352170 97094 352226
rect 97150 352170 97218 352226
rect 97274 352170 97342 352226
rect 97398 352170 97494 352226
rect 96874 352102 97494 352170
rect 96874 352046 96970 352102
rect 97026 352046 97094 352102
rect 97150 352046 97218 352102
rect 97274 352046 97342 352102
rect 97398 352046 97494 352102
rect 96874 351978 97494 352046
rect 96874 351922 96970 351978
rect 97026 351922 97094 351978
rect 97150 351922 97218 351978
rect 97274 351922 97342 351978
rect 97398 351922 97494 351978
rect 96874 334350 97494 351922
rect 100528 352350 100848 352384
rect 100528 352294 100598 352350
rect 100654 352294 100722 352350
rect 100778 352294 100848 352350
rect 100528 352226 100848 352294
rect 100528 352170 100598 352226
rect 100654 352170 100722 352226
rect 100778 352170 100848 352226
rect 100528 352102 100848 352170
rect 100528 352046 100598 352102
rect 100654 352046 100722 352102
rect 100778 352046 100848 352102
rect 100528 351978 100848 352046
rect 100528 351922 100598 351978
rect 100654 351922 100722 351978
rect 100778 351922 100848 351978
rect 100528 351888 100848 351922
rect 111154 346350 111774 363922
rect 115888 364350 116208 364384
rect 115888 364294 115958 364350
rect 116014 364294 116082 364350
rect 116138 364294 116208 364350
rect 115888 364226 116208 364294
rect 115888 364170 115958 364226
rect 116014 364170 116082 364226
rect 116138 364170 116208 364226
rect 115888 364102 116208 364170
rect 115888 364046 115958 364102
rect 116014 364046 116082 364102
rect 116138 364046 116208 364102
rect 115888 363978 116208 364046
rect 115888 363922 115958 363978
rect 116014 363922 116082 363978
rect 116138 363922 116208 363978
rect 115888 363888 116208 363922
rect 146608 364350 146928 364384
rect 146608 364294 146678 364350
rect 146734 364294 146802 364350
rect 146858 364294 146928 364350
rect 146608 364226 146928 364294
rect 146608 364170 146678 364226
rect 146734 364170 146802 364226
rect 146858 364170 146928 364226
rect 146608 364102 146928 364170
rect 146608 364046 146678 364102
rect 146734 364046 146802 364102
rect 146858 364046 146928 364102
rect 146608 363978 146928 364046
rect 146608 363922 146678 363978
rect 146734 363922 146802 363978
rect 146858 363922 146928 363978
rect 146608 363888 146928 363922
rect 177328 364350 177648 364384
rect 177328 364294 177398 364350
rect 177454 364294 177522 364350
rect 177578 364294 177648 364350
rect 177328 364226 177648 364294
rect 177328 364170 177398 364226
rect 177454 364170 177522 364226
rect 177578 364170 177648 364226
rect 177328 364102 177648 364170
rect 177328 364046 177398 364102
rect 177454 364046 177522 364102
rect 177578 364046 177648 364102
rect 177328 363978 177648 364046
rect 177328 363922 177398 363978
rect 177454 363922 177522 363978
rect 177578 363922 177648 363978
rect 177328 363888 177648 363922
rect 208048 364350 208368 364384
rect 208048 364294 208118 364350
rect 208174 364294 208242 364350
rect 208298 364294 208368 364350
rect 208048 364226 208368 364294
rect 208048 364170 208118 364226
rect 208174 364170 208242 364226
rect 208298 364170 208368 364226
rect 208048 364102 208368 364170
rect 208048 364046 208118 364102
rect 208174 364046 208242 364102
rect 208298 364046 208368 364102
rect 208048 363978 208368 364046
rect 208048 363922 208118 363978
rect 208174 363922 208242 363978
rect 208298 363922 208368 363978
rect 208048 363888 208368 363922
rect 238768 364350 239088 364384
rect 238768 364294 238838 364350
rect 238894 364294 238962 364350
rect 239018 364294 239088 364350
rect 238768 364226 239088 364294
rect 238768 364170 238838 364226
rect 238894 364170 238962 364226
rect 239018 364170 239088 364226
rect 238768 364102 239088 364170
rect 238768 364046 238838 364102
rect 238894 364046 238962 364102
rect 239018 364046 239088 364102
rect 238768 363978 239088 364046
rect 238768 363922 238838 363978
rect 238894 363922 238962 363978
rect 239018 363922 239088 363978
rect 238768 363888 239088 363922
rect 269488 364350 269808 364384
rect 269488 364294 269558 364350
rect 269614 364294 269682 364350
rect 269738 364294 269808 364350
rect 269488 364226 269808 364294
rect 269488 364170 269558 364226
rect 269614 364170 269682 364226
rect 269738 364170 269808 364226
rect 269488 364102 269808 364170
rect 269488 364046 269558 364102
rect 269614 364046 269682 364102
rect 269738 364046 269808 364102
rect 269488 363978 269808 364046
rect 269488 363922 269558 363978
rect 269614 363922 269682 363978
rect 269738 363922 269808 363978
rect 269488 363888 269808 363922
rect 300208 364350 300528 364384
rect 300208 364294 300278 364350
rect 300334 364294 300402 364350
rect 300458 364294 300528 364350
rect 300208 364226 300528 364294
rect 300208 364170 300278 364226
rect 300334 364170 300402 364226
rect 300458 364170 300528 364226
rect 300208 364102 300528 364170
rect 300208 364046 300278 364102
rect 300334 364046 300402 364102
rect 300458 364046 300528 364102
rect 300208 363978 300528 364046
rect 300208 363922 300278 363978
rect 300334 363922 300402 363978
rect 300458 363922 300528 363978
rect 300208 363888 300528 363922
rect 330928 364350 331248 364384
rect 330928 364294 330998 364350
rect 331054 364294 331122 364350
rect 331178 364294 331248 364350
rect 330928 364226 331248 364294
rect 330928 364170 330998 364226
rect 331054 364170 331122 364226
rect 331178 364170 331248 364226
rect 330928 364102 331248 364170
rect 330928 364046 330998 364102
rect 331054 364046 331122 364102
rect 331178 364046 331248 364102
rect 330928 363978 331248 364046
rect 330928 363922 330998 363978
rect 331054 363922 331122 363978
rect 331178 363922 331248 363978
rect 330928 363888 331248 363922
rect 361648 364350 361968 364384
rect 361648 364294 361718 364350
rect 361774 364294 361842 364350
rect 361898 364294 361968 364350
rect 361648 364226 361968 364294
rect 361648 364170 361718 364226
rect 361774 364170 361842 364226
rect 361898 364170 361968 364226
rect 361648 364102 361968 364170
rect 361648 364046 361718 364102
rect 361774 364046 361842 364102
rect 361898 364046 361968 364102
rect 361648 363978 361968 364046
rect 361648 363922 361718 363978
rect 361774 363922 361842 363978
rect 361898 363922 361968 363978
rect 361648 363888 361968 363922
rect 392368 364350 392688 364384
rect 392368 364294 392438 364350
rect 392494 364294 392562 364350
rect 392618 364294 392688 364350
rect 392368 364226 392688 364294
rect 392368 364170 392438 364226
rect 392494 364170 392562 364226
rect 392618 364170 392688 364226
rect 392368 364102 392688 364170
rect 392368 364046 392438 364102
rect 392494 364046 392562 364102
rect 392618 364046 392688 364102
rect 392368 363978 392688 364046
rect 392368 363922 392438 363978
rect 392494 363922 392562 363978
rect 392618 363922 392688 363978
rect 392368 363888 392688 363922
rect 423088 364350 423408 364384
rect 423088 364294 423158 364350
rect 423214 364294 423282 364350
rect 423338 364294 423408 364350
rect 423088 364226 423408 364294
rect 423088 364170 423158 364226
rect 423214 364170 423282 364226
rect 423338 364170 423408 364226
rect 423088 364102 423408 364170
rect 423088 364046 423158 364102
rect 423214 364046 423282 364102
rect 423338 364046 423408 364102
rect 423088 363978 423408 364046
rect 423088 363922 423158 363978
rect 423214 363922 423282 363978
rect 423338 363922 423408 363978
rect 423088 363888 423408 363922
rect 453808 364350 454128 364384
rect 453808 364294 453878 364350
rect 453934 364294 454002 364350
rect 454058 364294 454128 364350
rect 453808 364226 454128 364294
rect 453808 364170 453878 364226
rect 453934 364170 454002 364226
rect 454058 364170 454128 364226
rect 453808 364102 454128 364170
rect 453808 364046 453878 364102
rect 453934 364046 454002 364102
rect 454058 364046 454128 364102
rect 453808 363978 454128 364046
rect 453808 363922 453878 363978
rect 453934 363922 454002 363978
rect 454058 363922 454128 363978
rect 453808 363888 454128 363922
rect 484528 364350 484848 364384
rect 484528 364294 484598 364350
rect 484654 364294 484722 364350
rect 484778 364294 484848 364350
rect 484528 364226 484848 364294
rect 484528 364170 484598 364226
rect 484654 364170 484722 364226
rect 484778 364170 484848 364226
rect 484528 364102 484848 364170
rect 484528 364046 484598 364102
rect 484654 364046 484722 364102
rect 484778 364046 484848 364102
rect 484528 363978 484848 364046
rect 484528 363922 484598 363978
rect 484654 363922 484722 363978
rect 484778 363922 484848 363978
rect 484528 363888 484848 363922
rect 515248 364350 515568 364384
rect 515248 364294 515318 364350
rect 515374 364294 515442 364350
rect 515498 364294 515568 364350
rect 515248 364226 515568 364294
rect 515248 364170 515318 364226
rect 515374 364170 515442 364226
rect 515498 364170 515568 364226
rect 515248 364102 515568 364170
rect 515248 364046 515318 364102
rect 515374 364046 515442 364102
rect 515498 364046 515568 364102
rect 515248 363978 515568 364046
rect 515248 363922 515318 363978
rect 515374 363922 515442 363978
rect 515498 363922 515568 363978
rect 515248 363888 515568 363922
rect 545968 364350 546288 364384
rect 545968 364294 546038 364350
rect 546094 364294 546162 364350
rect 546218 364294 546288 364350
rect 545968 364226 546288 364294
rect 545968 364170 546038 364226
rect 546094 364170 546162 364226
rect 546218 364170 546288 364226
rect 545968 364102 546288 364170
rect 545968 364046 546038 364102
rect 546094 364046 546162 364102
rect 546218 364046 546288 364102
rect 545968 363978 546288 364046
rect 545968 363922 546038 363978
rect 546094 363922 546162 363978
rect 546218 363922 546288 363978
rect 545968 363888 546288 363922
rect 561154 364350 561774 381922
rect 561154 364294 561250 364350
rect 561306 364294 561374 364350
rect 561430 364294 561498 364350
rect 561554 364294 561622 364350
rect 561678 364294 561774 364350
rect 561154 364226 561774 364294
rect 561154 364170 561250 364226
rect 561306 364170 561374 364226
rect 561430 364170 561498 364226
rect 561554 364170 561622 364226
rect 561678 364170 561774 364226
rect 561154 364102 561774 364170
rect 561154 364046 561250 364102
rect 561306 364046 561374 364102
rect 561430 364046 561498 364102
rect 561554 364046 561622 364102
rect 561678 364046 561774 364102
rect 561154 363978 561774 364046
rect 561154 363922 561250 363978
rect 561306 363922 561374 363978
rect 561430 363922 561498 363978
rect 561554 363922 561622 363978
rect 561678 363922 561774 363978
rect 131248 352350 131568 352384
rect 131248 352294 131318 352350
rect 131374 352294 131442 352350
rect 131498 352294 131568 352350
rect 131248 352226 131568 352294
rect 131248 352170 131318 352226
rect 131374 352170 131442 352226
rect 131498 352170 131568 352226
rect 131248 352102 131568 352170
rect 131248 352046 131318 352102
rect 131374 352046 131442 352102
rect 131498 352046 131568 352102
rect 131248 351978 131568 352046
rect 131248 351922 131318 351978
rect 131374 351922 131442 351978
rect 131498 351922 131568 351978
rect 131248 351888 131568 351922
rect 161968 352350 162288 352384
rect 161968 352294 162038 352350
rect 162094 352294 162162 352350
rect 162218 352294 162288 352350
rect 161968 352226 162288 352294
rect 161968 352170 162038 352226
rect 162094 352170 162162 352226
rect 162218 352170 162288 352226
rect 161968 352102 162288 352170
rect 161968 352046 162038 352102
rect 162094 352046 162162 352102
rect 162218 352046 162288 352102
rect 161968 351978 162288 352046
rect 161968 351922 162038 351978
rect 162094 351922 162162 351978
rect 162218 351922 162288 351978
rect 161968 351888 162288 351922
rect 192688 352350 193008 352384
rect 192688 352294 192758 352350
rect 192814 352294 192882 352350
rect 192938 352294 193008 352350
rect 192688 352226 193008 352294
rect 192688 352170 192758 352226
rect 192814 352170 192882 352226
rect 192938 352170 193008 352226
rect 192688 352102 193008 352170
rect 192688 352046 192758 352102
rect 192814 352046 192882 352102
rect 192938 352046 193008 352102
rect 192688 351978 193008 352046
rect 192688 351922 192758 351978
rect 192814 351922 192882 351978
rect 192938 351922 193008 351978
rect 192688 351888 193008 351922
rect 223408 352350 223728 352384
rect 223408 352294 223478 352350
rect 223534 352294 223602 352350
rect 223658 352294 223728 352350
rect 223408 352226 223728 352294
rect 223408 352170 223478 352226
rect 223534 352170 223602 352226
rect 223658 352170 223728 352226
rect 223408 352102 223728 352170
rect 223408 352046 223478 352102
rect 223534 352046 223602 352102
rect 223658 352046 223728 352102
rect 223408 351978 223728 352046
rect 223408 351922 223478 351978
rect 223534 351922 223602 351978
rect 223658 351922 223728 351978
rect 223408 351888 223728 351922
rect 254128 352350 254448 352384
rect 254128 352294 254198 352350
rect 254254 352294 254322 352350
rect 254378 352294 254448 352350
rect 254128 352226 254448 352294
rect 254128 352170 254198 352226
rect 254254 352170 254322 352226
rect 254378 352170 254448 352226
rect 254128 352102 254448 352170
rect 254128 352046 254198 352102
rect 254254 352046 254322 352102
rect 254378 352046 254448 352102
rect 254128 351978 254448 352046
rect 254128 351922 254198 351978
rect 254254 351922 254322 351978
rect 254378 351922 254448 351978
rect 254128 351888 254448 351922
rect 284848 352350 285168 352384
rect 284848 352294 284918 352350
rect 284974 352294 285042 352350
rect 285098 352294 285168 352350
rect 284848 352226 285168 352294
rect 284848 352170 284918 352226
rect 284974 352170 285042 352226
rect 285098 352170 285168 352226
rect 284848 352102 285168 352170
rect 284848 352046 284918 352102
rect 284974 352046 285042 352102
rect 285098 352046 285168 352102
rect 284848 351978 285168 352046
rect 284848 351922 284918 351978
rect 284974 351922 285042 351978
rect 285098 351922 285168 351978
rect 284848 351888 285168 351922
rect 315568 352350 315888 352384
rect 315568 352294 315638 352350
rect 315694 352294 315762 352350
rect 315818 352294 315888 352350
rect 315568 352226 315888 352294
rect 315568 352170 315638 352226
rect 315694 352170 315762 352226
rect 315818 352170 315888 352226
rect 315568 352102 315888 352170
rect 315568 352046 315638 352102
rect 315694 352046 315762 352102
rect 315818 352046 315888 352102
rect 315568 351978 315888 352046
rect 315568 351922 315638 351978
rect 315694 351922 315762 351978
rect 315818 351922 315888 351978
rect 315568 351888 315888 351922
rect 346288 352350 346608 352384
rect 346288 352294 346358 352350
rect 346414 352294 346482 352350
rect 346538 352294 346608 352350
rect 346288 352226 346608 352294
rect 346288 352170 346358 352226
rect 346414 352170 346482 352226
rect 346538 352170 346608 352226
rect 346288 352102 346608 352170
rect 346288 352046 346358 352102
rect 346414 352046 346482 352102
rect 346538 352046 346608 352102
rect 346288 351978 346608 352046
rect 346288 351922 346358 351978
rect 346414 351922 346482 351978
rect 346538 351922 346608 351978
rect 346288 351888 346608 351922
rect 377008 352350 377328 352384
rect 377008 352294 377078 352350
rect 377134 352294 377202 352350
rect 377258 352294 377328 352350
rect 377008 352226 377328 352294
rect 377008 352170 377078 352226
rect 377134 352170 377202 352226
rect 377258 352170 377328 352226
rect 377008 352102 377328 352170
rect 377008 352046 377078 352102
rect 377134 352046 377202 352102
rect 377258 352046 377328 352102
rect 377008 351978 377328 352046
rect 377008 351922 377078 351978
rect 377134 351922 377202 351978
rect 377258 351922 377328 351978
rect 377008 351888 377328 351922
rect 407728 352350 408048 352384
rect 407728 352294 407798 352350
rect 407854 352294 407922 352350
rect 407978 352294 408048 352350
rect 407728 352226 408048 352294
rect 407728 352170 407798 352226
rect 407854 352170 407922 352226
rect 407978 352170 408048 352226
rect 407728 352102 408048 352170
rect 407728 352046 407798 352102
rect 407854 352046 407922 352102
rect 407978 352046 408048 352102
rect 407728 351978 408048 352046
rect 407728 351922 407798 351978
rect 407854 351922 407922 351978
rect 407978 351922 408048 351978
rect 407728 351888 408048 351922
rect 438448 352350 438768 352384
rect 438448 352294 438518 352350
rect 438574 352294 438642 352350
rect 438698 352294 438768 352350
rect 438448 352226 438768 352294
rect 438448 352170 438518 352226
rect 438574 352170 438642 352226
rect 438698 352170 438768 352226
rect 438448 352102 438768 352170
rect 438448 352046 438518 352102
rect 438574 352046 438642 352102
rect 438698 352046 438768 352102
rect 438448 351978 438768 352046
rect 438448 351922 438518 351978
rect 438574 351922 438642 351978
rect 438698 351922 438768 351978
rect 438448 351888 438768 351922
rect 469168 352350 469488 352384
rect 469168 352294 469238 352350
rect 469294 352294 469362 352350
rect 469418 352294 469488 352350
rect 469168 352226 469488 352294
rect 469168 352170 469238 352226
rect 469294 352170 469362 352226
rect 469418 352170 469488 352226
rect 469168 352102 469488 352170
rect 469168 352046 469238 352102
rect 469294 352046 469362 352102
rect 469418 352046 469488 352102
rect 469168 351978 469488 352046
rect 469168 351922 469238 351978
rect 469294 351922 469362 351978
rect 469418 351922 469488 351978
rect 469168 351888 469488 351922
rect 499888 352350 500208 352384
rect 499888 352294 499958 352350
rect 500014 352294 500082 352350
rect 500138 352294 500208 352350
rect 499888 352226 500208 352294
rect 499888 352170 499958 352226
rect 500014 352170 500082 352226
rect 500138 352170 500208 352226
rect 499888 352102 500208 352170
rect 499888 352046 499958 352102
rect 500014 352046 500082 352102
rect 500138 352046 500208 352102
rect 499888 351978 500208 352046
rect 499888 351922 499958 351978
rect 500014 351922 500082 351978
rect 500138 351922 500208 351978
rect 499888 351888 500208 351922
rect 530608 352350 530928 352384
rect 530608 352294 530678 352350
rect 530734 352294 530802 352350
rect 530858 352294 530928 352350
rect 530608 352226 530928 352294
rect 530608 352170 530678 352226
rect 530734 352170 530802 352226
rect 530858 352170 530928 352226
rect 530608 352102 530928 352170
rect 530608 352046 530678 352102
rect 530734 352046 530802 352102
rect 530858 352046 530928 352102
rect 530608 351978 530928 352046
rect 530608 351922 530678 351978
rect 530734 351922 530802 351978
rect 530858 351922 530928 351978
rect 530608 351888 530928 351922
rect 111154 346294 111250 346350
rect 111306 346294 111374 346350
rect 111430 346294 111498 346350
rect 111554 346294 111622 346350
rect 111678 346294 111774 346350
rect 111154 346226 111774 346294
rect 111154 346170 111250 346226
rect 111306 346170 111374 346226
rect 111430 346170 111498 346226
rect 111554 346170 111622 346226
rect 111678 346170 111774 346226
rect 111154 346102 111774 346170
rect 111154 346046 111250 346102
rect 111306 346046 111374 346102
rect 111430 346046 111498 346102
rect 111554 346046 111622 346102
rect 111678 346046 111774 346102
rect 111154 345978 111774 346046
rect 111154 345922 111250 345978
rect 111306 345922 111374 345978
rect 111430 345922 111498 345978
rect 111554 345922 111622 345978
rect 111678 345922 111774 345978
rect 96874 334294 96970 334350
rect 97026 334294 97094 334350
rect 97150 334294 97218 334350
rect 97274 334294 97342 334350
rect 97398 334294 97494 334350
rect 96874 334226 97494 334294
rect 96874 334170 96970 334226
rect 97026 334170 97094 334226
rect 97150 334170 97218 334226
rect 97274 334170 97342 334226
rect 97398 334170 97494 334226
rect 96874 334102 97494 334170
rect 96874 334046 96970 334102
rect 97026 334046 97094 334102
rect 97150 334046 97218 334102
rect 97274 334046 97342 334102
rect 97398 334046 97494 334102
rect 96874 333978 97494 334046
rect 96874 333922 96970 333978
rect 97026 333922 97094 333978
rect 97150 333922 97218 333978
rect 97274 333922 97342 333978
rect 97398 333922 97494 333978
rect 96874 316350 97494 333922
rect 100528 334350 100848 334384
rect 100528 334294 100598 334350
rect 100654 334294 100722 334350
rect 100778 334294 100848 334350
rect 100528 334226 100848 334294
rect 100528 334170 100598 334226
rect 100654 334170 100722 334226
rect 100778 334170 100848 334226
rect 100528 334102 100848 334170
rect 100528 334046 100598 334102
rect 100654 334046 100722 334102
rect 100778 334046 100848 334102
rect 100528 333978 100848 334046
rect 100528 333922 100598 333978
rect 100654 333922 100722 333978
rect 100778 333922 100848 333978
rect 100528 333888 100848 333922
rect 111154 328350 111774 345922
rect 115888 346350 116208 346384
rect 115888 346294 115958 346350
rect 116014 346294 116082 346350
rect 116138 346294 116208 346350
rect 115888 346226 116208 346294
rect 115888 346170 115958 346226
rect 116014 346170 116082 346226
rect 116138 346170 116208 346226
rect 115888 346102 116208 346170
rect 115888 346046 115958 346102
rect 116014 346046 116082 346102
rect 116138 346046 116208 346102
rect 115888 345978 116208 346046
rect 115888 345922 115958 345978
rect 116014 345922 116082 345978
rect 116138 345922 116208 345978
rect 115888 345888 116208 345922
rect 146608 346350 146928 346384
rect 146608 346294 146678 346350
rect 146734 346294 146802 346350
rect 146858 346294 146928 346350
rect 146608 346226 146928 346294
rect 146608 346170 146678 346226
rect 146734 346170 146802 346226
rect 146858 346170 146928 346226
rect 146608 346102 146928 346170
rect 146608 346046 146678 346102
rect 146734 346046 146802 346102
rect 146858 346046 146928 346102
rect 146608 345978 146928 346046
rect 146608 345922 146678 345978
rect 146734 345922 146802 345978
rect 146858 345922 146928 345978
rect 146608 345888 146928 345922
rect 177328 346350 177648 346384
rect 177328 346294 177398 346350
rect 177454 346294 177522 346350
rect 177578 346294 177648 346350
rect 177328 346226 177648 346294
rect 177328 346170 177398 346226
rect 177454 346170 177522 346226
rect 177578 346170 177648 346226
rect 177328 346102 177648 346170
rect 177328 346046 177398 346102
rect 177454 346046 177522 346102
rect 177578 346046 177648 346102
rect 177328 345978 177648 346046
rect 177328 345922 177398 345978
rect 177454 345922 177522 345978
rect 177578 345922 177648 345978
rect 177328 345888 177648 345922
rect 208048 346350 208368 346384
rect 208048 346294 208118 346350
rect 208174 346294 208242 346350
rect 208298 346294 208368 346350
rect 208048 346226 208368 346294
rect 208048 346170 208118 346226
rect 208174 346170 208242 346226
rect 208298 346170 208368 346226
rect 208048 346102 208368 346170
rect 208048 346046 208118 346102
rect 208174 346046 208242 346102
rect 208298 346046 208368 346102
rect 208048 345978 208368 346046
rect 208048 345922 208118 345978
rect 208174 345922 208242 345978
rect 208298 345922 208368 345978
rect 208048 345888 208368 345922
rect 238768 346350 239088 346384
rect 238768 346294 238838 346350
rect 238894 346294 238962 346350
rect 239018 346294 239088 346350
rect 238768 346226 239088 346294
rect 238768 346170 238838 346226
rect 238894 346170 238962 346226
rect 239018 346170 239088 346226
rect 238768 346102 239088 346170
rect 238768 346046 238838 346102
rect 238894 346046 238962 346102
rect 239018 346046 239088 346102
rect 238768 345978 239088 346046
rect 238768 345922 238838 345978
rect 238894 345922 238962 345978
rect 239018 345922 239088 345978
rect 238768 345888 239088 345922
rect 269488 346350 269808 346384
rect 269488 346294 269558 346350
rect 269614 346294 269682 346350
rect 269738 346294 269808 346350
rect 269488 346226 269808 346294
rect 269488 346170 269558 346226
rect 269614 346170 269682 346226
rect 269738 346170 269808 346226
rect 269488 346102 269808 346170
rect 269488 346046 269558 346102
rect 269614 346046 269682 346102
rect 269738 346046 269808 346102
rect 269488 345978 269808 346046
rect 269488 345922 269558 345978
rect 269614 345922 269682 345978
rect 269738 345922 269808 345978
rect 269488 345888 269808 345922
rect 300208 346350 300528 346384
rect 300208 346294 300278 346350
rect 300334 346294 300402 346350
rect 300458 346294 300528 346350
rect 300208 346226 300528 346294
rect 300208 346170 300278 346226
rect 300334 346170 300402 346226
rect 300458 346170 300528 346226
rect 300208 346102 300528 346170
rect 300208 346046 300278 346102
rect 300334 346046 300402 346102
rect 300458 346046 300528 346102
rect 300208 345978 300528 346046
rect 300208 345922 300278 345978
rect 300334 345922 300402 345978
rect 300458 345922 300528 345978
rect 300208 345888 300528 345922
rect 330928 346350 331248 346384
rect 330928 346294 330998 346350
rect 331054 346294 331122 346350
rect 331178 346294 331248 346350
rect 330928 346226 331248 346294
rect 330928 346170 330998 346226
rect 331054 346170 331122 346226
rect 331178 346170 331248 346226
rect 330928 346102 331248 346170
rect 330928 346046 330998 346102
rect 331054 346046 331122 346102
rect 331178 346046 331248 346102
rect 330928 345978 331248 346046
rect 330928 345922 330998 345978
rect 331054 345922 331122 345978
rect 331178 345922 331248 345978
rect 330928 345888 331248 345922
rect 361648 346350 361968 346384
rect 361648 346294 361718 346350
rect 361774 346294 361842 346350
rect 361898 346294 361968 346350
rect 361648 346226 361968 346294
rect 361648 346170 361718 346226
rect 361774 346170 361842 346226
rect 361898 346170 361968 346226
rect 361648 346102 361968 346170
rect 361648 346046 361718 346102
rect 361774 346046 361842 346102
rect 361898 346046 361968 346102
rect 361648 345978 361968 346046
rect 361648 345922 361718 345978
rect 361774 345922 361842 345978
rect 361898 345922 361968 345978
rect 361648 345888 361968 345922
rect 392368 346350 392688 346384
rect 392368 346294 392438 346350
rect 392494 346294 392562 346350
rect 392618 346294 392688 346350
rect 392368 346226 392688 346294
rect 392368 346170 392438 346226
rect 392494 346170 392562 346226
rect 392618 346170 392688 346226
rect 392368 346102 392688 346170
rect 392368 346046 392438 346102
rect 392494 346046 392562 346102
rect 392618 346046 392688 346102
rect 392368 345978 392688 346046
rect 392368 345922 392438 345978
rect 392494 345922 392562 345978
rect 392618 345922 392688 345978
rect 392368 345888 392688 345922
rect 423088 346350 423408 346384
rect 423088 346294 423158 346350
rect 423214 346294 423282 346350
rect 423338 346294 423408 346350
rect 423088 346226 423408 346294
rect 423088 346170 423158 346226
rect 423214 346170 423282 346226
rect 423338 346170 423408 346226
rect 423088 346102 423408 346170
rect 423088 346046 423158 346102
rect 423214 346046 423282 346102
rect 423338 346046 423408 346102
rect 423088 345978 423408 346046
rect 423088 345922 423158 345978
rect 423214 345922 423282 345978
rect 423338 345922 423408 345978
rect 423088 345888 423408 345922
rect 453808 346350 454128 346384
rect 453808 346294 453878 346350
rect 453934 346294 454002 346350
rect 454058 346294 454128 346350
rect 453808 346226 454128 346294
rect 453808 346170 453878 346226
rect 453934 346170 454002 346226
rect 454058 346170 454128 346226
rect 453808 346102 454128 346170
rect 453808 346046 453878 346102
rect 453934 346046 454002 346102
rect 454058 346046 454128 346102
rect 453808 345978 454128 346046
rect 453808 345922 453878 345978
rect 453934 345922 454002 345978
rect 454058 345922 454128 345978
rect 453808 345888 454128 345922
rect 484528 346350 484848 346384
rect 484528 346294 484598 346350
rect 484654 346294 484722 346350
rect 484778 346294 484848 346350
rect 484528 346226 484848 346294
rect 484528 346170 484598 346226
rect 484654 346170 484722 346226
rect 484778 346170 484848 346226
rect 484528 346102 484848 346170
rect 484528 346046 484598 346102
rect 484654 346046 484722 346102
rect 484778 346046 484848 346102
rect 484528 345978 484848 346046
rect 484528 345922 484598 345978
rect 484654 345922 484722 345978
rect 484778 345922 484848 345978
rect 484528 345888 484848 345922
rect 515248 346350 515568 346384
rect 515248 346294 515318 346350
rect 515374 346294 515442 346350
rect 515498 346294 515568 346350
rect 515248 346226 515568 346294
rect 515248 346170 515318 346226
rect 515374 346170 515442 346226
rect 515498 346170 515568 346226
rect 515248 346102 515568 346170
rect 515248 346046 515318 346102
rect 515374 346046 515442 346102
rect 515498 346046 515568 346102
rect 515248 345978 515568 346046
rect 515248 345922 515318 345978
rect 515374 345922 515442 345978
rect 515498 345922 515568 345978
rect 515248 345888 515568 345922
rect 545968 346350 546288 346384
rect 545968 346294 546038 346350
rect 546094 346294 546162 346350
rect 546218 346294 546288 346350
rect 545968 346226 546288 346294
rect 545968 346170 546038 346226
rect 546094 346170 546162 346226
rect 546218 346170 546288 346226
rect 545968 346102 546288 346170
rect 545968 346046 546038 346102
rect 546094 346046 546162 346102
rect 546218 346046 546288 346102
rect 545968 345978 546288 346046
rect 545968 345922 546038 345978
rect 546094 345922 546162 345978
rect 546218 345922 546288 345978
rect 545968 345888 546288 345922
rect 561154 346350 561774 363922
rect 561154 346294 561250 346350
rect 561306 346294 561374 346350
rect 561430 346294 561498 346350
rect 561554 346294 561622 346350
rect 561678 346294 561774 346350
rect 561154 346226 561774 346294
rect 561154 346170 561250 346226
rect 561306 346170 561374 346226
rect 561430 346170 561498 346226
rect 561554 346170 561622 346226
rect 561678 346170 561774 346226
rect 561154 346102 561774 346170
rect 561154 346046 561250 346102
rect 561306 346046 561374 346102
rect 561430 346046 561498 346102
rect 561554 346046 561622 346102
rect 561678 346046 561774 346102
rect 561154 345978 561774 346046
rect 561154 345922 561250 345978
rect 561306 345922 561374 345978
rect 561430 345922 561498 345978
rect 561554 345922 561622 345978
rect 561678 345922 561774 345978
rect 131248 334350 131568 334384
rect 131248 334294 131318 334350
rect 131374 334294 131442 334350
rect 131498 334294 131568 334350
rect 131248 334226 131568 334294
rect 131248 334170 131318 334226
rect 131374 334170 131442 334226
rect 131498 334170 131568 334226
rect 131248 334102 131568 334170
rect 131248 334046 131318 334102
rect 131374 334046 131442 334102
rect 131498 334046 131568 334102
rect 131248 333978 131568 334046
rect 131248 333922 131318 333978
rect 131374 333922 131442 333978
rect 131498 333922 131568 333978
rect 131248 333888 131568 333922
rect 161968 334350 162288 334384
rect 161968 334294 162038 334350
rect 162094 334294 162162 334350
rect 162218 334294 162288 334350
rect 161968 334226 162288 334294
rect 161968 334170 162038 334226
rect 162094 334170 162162 334226
rect 162218 334170 162288 334226
rect 161968 334102 162288 334170
rect 161968 334046 162038 334102
rect 162094 334046 162162 334102
rect 162218 334046 162288 334102
rect 161968 333978 162288 334046
rect 161968 333922 162038 333978
rect 162094 333922 162162 333978
rect 162218 333922 162288 333978
rect 161968 333888 162288 333922
rect 192688 334350 193008 334384
rect 192688 334294 192758 334350
rect 192814 334294 192882 334350
rect 192938 334294 193008 334350
rect 192688 334226 193008 334294
rect 192688 334170 192758 334226
rect 192814 334170 192882 334226
rect 192938 334170 193008 334226
rect 192688 334102 193008 334170
rect 192688 334046 192758 334102
rect 192814 334046 192882 334102
rect 192938 334046 193008 334102
rect 192688 333978 193008 334046
rect 192688 333922 192758 333978
rect 192814 333922 192882 333978
rect 192938 333922 193008 333978
rect 192688 333888 193008 333922
rect 223408 334350 223728 334384
rect 223408 334294 223478 334350
rect 223534 334294 223602 334350
rect 223658 334294 223728 334350
rect 223408 334226 223728 334294
rect 223408 334170 223478 334226
rect 223534 334170 223602 334226
rect 223658 334170 223728 334226
rect 223408 334102 223728 334170
rect 223408 334046 223478 334102
rect 223534 334046 223602 334102
rect 223658 334046 223728 334102
rect 223408 333978 223728 334046
rect 223408 333922 223478 333978
rect 223534 333922 223602 333978
rect 223658 333922 223728 333978
rect 223408 333888 223728 333922
rect 254128 334350 254448 334384
rect 254128 334294 254198 334350
rect 254254 334294 254322 334350
rect 254378 334294 254448 334350
rect 254128 334226 254448 334294
rect 254128 334170 254198 334226
rect 254254 334170 254322 334226
rect 254378 334170 254448 334226
rect 254128 334102 254448 334170
rect 254128 334046 254198 334102
rect 254254 334046 254322 334102
rect 254378 334046 254448 334102
rect 254128 333978 254448 334046
rect 254128 333922 254198 333978
rect 254254 333922 254322 333978
rect 254378 333922 254448 333978
rect 254128 333888 254448 333922
rect 284848 334350 285168 334384
rect 284848 334294 284918 334350
rect 284974 334294 285042 334350
rect 285098 334294 285168 334350
rect 284848 334226 285168 334294
rect 284848 334170 284918 334226
rect 284974 334170 285042 334226
rect 285098 334170 285168 334226
rect 284848 334102 285168 334170
rect 284848 334046 284918 334102
rect 284974 334046 285042 334102
rect 285098 334046 285168 334102
rect 284848 333978 285168 334046
rect 284848 333922 284918 333978
rect 284974 333922 285042 333978
rect 285098 333922 285168 333978
rect 284848 333888 285168 333922
rect 315568 334350 315888 334384
rect 315568 334294 315638 334350
rect 315694 334294 315762 334350
rect 315818 334294 315888 334350
rect 315568 334226 315888 334294
rect 315568 334170 315638 334226
rect 315694 334170 315762 334226
rect 315818 334170 315888 334226
rect 315568 334102 315888 334170
rect 315568 334046 315638 334102
rect 315694 334046 315762 334102
rect 315818 334046 315888 334102
rect 315568 333978 315888 334046
rect 315568 333922 315638 333978
rect 315694 333922 315762 333978
rect 315818 333922 315888 333978
rect 315568 333888 315888 333922
rect 346288 334350 346608 334384
rect 346288 334294 346358 334350
rect 346414 334294 346482 334350
rect 346538 334294 346608 334350
rect 346288 334226 346608 334294
rect 346288 334170 346358 334226
rect 346414 334170 346482 334226
rect 346538 334170 346608 334226
rect 346288 334102 346608 334170
rect 346288 334046 346358 334102
rect 346414 334046 346482 334102
rect 346538 334046 346608 334102
rect 346288 333978 346608 334046
rect 346288 333922 346358 333978
rect 346414 333922 346482 333978
rect 346538 333922 346608 333978
rect 346288 333888 346608 333922
rect 377008 334350 377328 334384
rect 377008 334294 377078 334350
rect 377134 334294 377202 334350
rect 377258 334294 377328 334350
rect 377008 334226 377328 334294
rect 377008 334170 377078 334226
rect 377134 334170 377202 334226
rect 377258 334170 377328 334226
rect 377008 334102 377328 334170
rect 377008 334046 377078 334102
rect 377134 334046 377202 334102
rect 377258 334046 377328 334102
rect 377008 333978 377328 334046
rect 377008 333922 377078 333978
rect 377134 333922 377202 333978
rect 377258 333922 377328 333978
rect 377008 333888 377328 333922
rect 407728 334350 408048 334384
rect 407728 334294 407798 334350
rect 407854 334294 407922 334350
rect 407978 334294 408048 334350
rect 407728 334226 408048 334294
rect 407728 334170 407798 334226
rect 407854 334170 407922 334226
rect 407978 334170 408048 334226
rect 407728 334102 408048 334170
rect 407728 334046 407798 334102
rect 407854 334046 407922 334102
rect 407978 334046 408048 334102
rect 407728 333978 408048 334046
rect 407728 333922 407798 333978
rect 407854 333922 407922 333978
rect 407978 333922 408048 333978
rect 407728 333888 408048 333922
rect 438448 334350 438768 334384
rect 438448 334294 438518 334350
rect 438574 334294 438642 334350
rect 438698 334294 438768 334350
rect 438448 334226 438768 334294
rect 438448 334170 438518 334226
rect 438574 334170 438642 334226
rect 438698 334170 438768 334226
rect 438448 334102 438768 334170
rect 438448 334046 438518 334102
rect 438574 334046 438642 334102
rect 438698 334046 438768 334102
rect 438448 333978 438768 334046
rect 438448 333922 438518 333978
rect 438574 333922 438642 333978
rect 438698 333922 438768 333978
rect 438448 333888 438768 333922
rect 469168 334350 469488 334384
rect 469168 334294 469238 334350
rect 469294 334294 469362 334350
rect 469418 334294 469488 334350
rect 469168 334226 469488 334294
rect 469168 334170 469238 334226
rect 469294 334170 469362 334226
rect 469418 334170 469488 334226
rect 469168 334102 469488 334170
rect 469168 334046 469238 334102
rect 469294 334046 469362 334102
rect 469418 334046 469488 334102
rect 469168 333978 469488 334046
rect 469168 333922 469238 333978
rect 469294 333922 469362 333978
rect 469418 333922 469488 333978
rect 469168 333888 469488 333922
rect 499888 334350 500208 334384
rect 499888 334294 499958 334350
rect 500014 334294 500082 334350
rect 500138 334294 500208 334350
rect 499888 334226 500208 334294
rect 499888 334170 499958 334226
rect 500014 334170 500082 334226
rect 500138 334170 500208 334226
rect 499888 334102 500208 334170
rect 499888 334046 499958 334102
rect 500014 334046 500082 334102
rect 500138 334046 500208 334102
rect 499888 333978 500208 334046
rect 499888 333922 499958 333978
rect 500014 333922 500082 333978
rect 500138 333922 500208 333978
rect 499888 333888 500208 333922
rect 530608 334350 530928 334384
rect 530608 334294 530678 334350
rect 530734 334294 530802 334350
rect 530858 334294 530928 334350
rect 530608 334226 530928 334294
rect 530608 334170 530678 334226
rect 530734 334170 530802 334226
rect 530858 334170 530928 334226
rect 530608 334102 530928 334170
rect 530608 334046 530678 334102
rect 530734 334046 530802 334102
rect 530858 334046 530928 334102
rect 530608 333978 530928 334046
rect 530608 333922 530678 333978
rect 530734 333922 530802 333978
rect 530858 333922 530928 333978
rect 530608 333888 530928 333922
rect 111154 328294 111250 328350
rect 111306 328294 111374 328350
rect 111430 328294 111498 328350
rect 111554 328294 111622 328350
rect 111678 328294 111774 328350
rect 111154 328226 111774 328294
rect 111154 328170 111250 328226
rect 111306 328170 111374 328226
rect 111430 328170 111498 328226
rect 111554 328170 111622 328226
rect 111678 328170 111774 328226
rect 111154 328102 111774 328170
rect 111154 328046 111250 328102
rect 111306 328046 111374 328102
rect 111430 328046 111498 328102
rect 111554 328046 111622 328102
rect 111678 328046 111774 328102
rect 111154 327978 111774 328046
rect 111154 327922 111250 327978
rect 111306 327922 111374 327978
rect 111430 327922 111498 327978
rect 111554 327922 111622 327978
rect 111678 327922 111774 327978
rect 96874 316294 96970 316350
rect 97026 316294 97094 316350
rect 97150 316294 97218 316350
rect 97274 316294 97342 316350
rect 97398 316294 97494 316350
rect 96874 316226 97494 316294
rect 96874 316170 96970 316226
rect 97026 316170 97094 316226
rect 97150 316170 97218 316226
rect 97274 316170 97342 316226
rect 97398 316170 97494 316226
rect 96874 316102 97494 316170
rect 96874 316046 96970 316102
rect 97026 316046 97094 316102
rect 97150 316046 97218 316102
rect 97274 316046 97342 316102
rect 97398 316046 97494 316102
rect 96874 315978 97494 316046
rect 96874 315922 96970 315978
rect 97026 315922 97094 315978
rect 97150 315922 97218 315978
rect 97274 315922 97342 315978
rect 97398 315922 97494 315978
rect 96874 298350 97494 315922
rect 100528 316350 100848 316384
rect 100528 316294 100598 316350
rect 100654 316294 100722 316350
rect 100778 316294 100848 316350
rect 100528 316226 100848 316294
rect 100528 316170 100598 316226
rect 100654 316170 100722 316226
rect 100778 316170 100848 316226
rect 100528 316102 100848 316170
rect 100528 316046 100598 316102
rect 100654 316046 100722 316102
rect 100778 316046 100848 316102
rect 100528 315978 100848 316046
rect 100528 315922 100598 315978
rect 100654 315922 100722 315978
rect 100778 315922 100848 315978
rect 100528 315888 100848 315922
rect 111154 310350 111774 327922
rect 115888 328350 116208 328384
rect 115888 328294 115958 328350
rect 116014 328294 116082 328350
rect 116138 328294 116208 328350
rect 115888 328226 116208 328294
rect 115888 328170 115958 328226
rect 116014 328170 116082 328226
rect 116138 328170 116208 328226
rect 115888 328102 116208 328170
rect 115888 328046 115958 328102
rect 116014 328046 116082 328102
rect 116138 328046 116208 328102
rect 115888 327978 116208 328046
rect 115888 327922 115958 327978
rect 116014 327922 116082 327978
rect 116138 327922 116208 327978
rect 115888 327888 116208 327922
rect 146608 328350 146928 328384
rect 146608 328294 146678 328350
rect 146734 328294 146802 328350
rect 146858 328294 146928 328350
rect 146608 328226 146928 328294
rect 146608 328170 146678 328226
rect 146734 328170 146802 328226
rect 146858 328170 146928 328226
rect 146608 328102 146928 328170
rect 146608 328046 146678 328102
rect 146734 328046 146802 328102
rect 146858 328046 146928 328102
rect 146608 327978 146928 328046
rect 146608 327922 146678 327978
rect 146734 327922 146802 327978
rect 146858 327922 146928 327978
rect 146608 327888 146928 327922
rect 177328 328350 177648 328384
rect 177328 328294 177398 328350
rect 177454 328294 177522 328350
rect 177578 328294 177648 328350
rect 177328 328226 177648 328294
rect 177328 328170 177398 328226
rect 177454 328170 177522 328226
rect 177578 328170 177648 328226
rect 177328 328102 177648 328170
rect 177328 328046 177398 328102
rect 177454 328046 177522 328102
rect 177578 328046 177648 328102
rect 177328 327978 177648 328046
rect 177328 327922 177398 327978
rect 177454 327922 177522 327978
rect 177578 327922 177648 327978
rect 177328 327888 177648 327922
rect 208048 328350 208368 328384
rect 208048 328294 208118 328350
rect 208174 328294 208242 328350
rect 208298 328294 208368 328350
rect 208048 328226 208368 328294
rect 208048 328170 208118 328226
rect 208174 328170 208242 328226
rect 208298 328170 208368 328226
rect 208048 328102 208368 328170
rect 208048 328046 208118 328102
rect 208174 328046 208242 328102
rect 208298 328046 208368 328102
rect 208048 327978 208368 328046
rect 208048 327922 208118 327978
rect 208174 327922 208242 327978
rect 208298 327922 208368 327978
rect 208048 327888 208368 327922
rect 238768 328350 239088 328384
rect 238768 328294 238838 328350
rect 238894 328294 238962 328350
rect 239018 328294 239088 328350
rect 238768 328226 239088 328294
rect 238768 328170 238838 328226
rect 238894 328170 238962 328226
rect 239018 328170 239088 328226
rect 238768 328102 239088 328170
rect 238768 328046 238838 328102
rect 238894 328046 238962 328102
rect 239018 328046 239088 328102
rect 238768 327978 239088 328046
rect 238768 327922 238838 327978
rect 238894 327922 238962 327978
rect 239018 327922 239088 327978
rect 238768 327888 239088 327922
rect 269488 328350 269808 328384
rect 269488 328294 269558 328350
rect 269614 328294 269682 328350
rect 269738 328294 269808 328350
rect 269488 328226 269808 328294
rect 269488 328170 269558 328226
rect 269614 328170 269682 328226
rect 269738 328170 269808 328226
rect 269488 328102 269808 328170
rect 269488 328046 269558 328102
rect 269614 328046 269682 328102
rect 269738 328046 269808 328102
rect 269488 327978 269808 328046
rect 269488 327922 269558 327978
rect 269614 327922 269682 327978
rect 269738 327922 269808 327978
rect 269488 327888 269808 327922
rect 300208 328350 300528 328384
rect 300208 328294 300278 328350
rect 300334 328294 300402 328350
rect 300458 328294 300528 328350
rect 300208 328226 300528 328294
rect 300208 328170 300278 328226
rect 300334 328170 300402 328226
rect 300458 328170 300528 328226
rect 300208 328102 300528 328170
rect 300208 328046 300278 328102
rect 300334 328046 300402 328102
rect 300458 328046 300528 328102
rect 300208 327978 300528 328046
rect 300208 327922 300278 327978
rect 300334 327922 300402 327978
rect 300458 327922 300528 327978
rect 300208 327888 300528 327922
rect 330928 328350 331248 328384
rect 330928 328294 330998 328350
rect 331054 328294 331122 328350
rect 331178 328294 331248 328350
rect 330928 328226 331248 328294
rect 330928 328170 330998 328226
rect 331054 328170 331122 328226
rect 331178 328170 331248 328226
rect 330928 328102 331248 328170
rect 330928 328046 330998 328102
rect 331054 328046 331122 328102
rect 331178 328046 331248 328102
rect 330928 327978 331248 328046
rect 330928 327922 330998 327978
rect 331054 327922 331122 327978
rect 331178 327922 331248 327978
rect 330928 327888 331248 327922
rect 361648 328350 361968 328384
rect 361648 328294 361718 328350
rect 361774 328294 361842 328350
rect 361898 328294 361968 328350
rect 361648 328226 361968 328294
rect 361648 328170 361718 328226
rect 361774 328170 361842 328226
rect 361898 328170 361968 328226
rect 361648 328102 361968 328170
rect 361648 328046 361718 328102
rect 361774 328046 361842 328102
rect 361898 328046 361968 328102
rect 361648 327978 361968 328046
rect 361648 327922 361718 327978
rect 361774 327922 361842 327978
rect 361898 327922 361968 327978
rect 361648 327888 361968 327922
rect 392368 328350 392688 328384
rect 392368 328294 392438 328350
rect 392494 328294 392562 328350
rect 392618 328294 392688 328350
rect 392368 328226 392688 328294
rect 392368 328170 392438 328226
rect 392494 328170 392562 328226
rect 392618 328170 392688 328226
rect 392368 328102 392688 328170
rect 392368 328046 392438 328102
rect 392494 328046 392562 328102
rect 392618 328046 392688 328102
rect 392368 327978 392688 328046
rect 392368 327922 392438 327978
rect 392494 327922 392562 327978
rect 392618 327922 392688 327978
rect 392368 327888 392688 327922
rect 423088 328350 423408 328384
rect 423088 328294 423158 328350
rect 423214 328294 423282 328350
rect 423338 328294 423408 328350
rect 423088 328226 423408 328294
rect 423088 328170 423158 328226
rect 423214 328170 423282 328226
rect 423338 328170 423408 328226
rect 423088 328102 423408 328170
rect 423088 328046 423158 328102
rect 423214 328046 423282 328102
rect 423338 328046 423408 328102
rect 423088 327978 423408 328046
rect 423088 327922 423158 327978
rect 423214 327922 423282 327978
rect 423338 327922 423408 327978
rect 423088 327888 423408 327922
rect 453808 328350 454128 328384
rect 453808 328294 453878 328350
rect 453934 328294 454002 328350
rect 454058 328294 454128 328350
rect 453808 328226 454128 328294
rect 453808 328170 453878 328226
rect 453934 328170 454002 328226
rect 454058 328170 454128 328226
rect 453808 328102 454128 328170
rect 453808 328046 453878 328102
rect 453934 328046 454002 328102
rect 454058 328046 454128 328102
rect 453808 327978 454128 328046
rect 453808 327922 453878 327978
rect 453934 327922 454002 327978
rect 454058 327922 454128 327978
rect 453808 327888 454128 327922
rect 484528 328350 484848 328384
rect 484528 328294 484598 328350
rect 484654 328294 484722 328350
rect 484778 328294 484848 328350
rect 484528 328226 484848 328294
rect 484528 328170 484598 328226
rect 484654 328170 484722 328226
rect 484778 328170 484848 328226
rect 484528 328102 484848 328170
rect 484528 328046 484598 328102
rect 484654 328046 484722 328102
rect 484778 328046 484848 328102
rect 484528 327978 484848 328046
rect 484528 327922 484598 327978
rect 484654 327922 484722 327978
rect 484778 327922 484848 327978
rect 484528 327888 484848 327922
rect 515248 328350 515568 328384
rect 515248 328294 515318 328350
rect 515374 328294 515442 328350
rect 515498 328294 515568 328350
rect 515248 328226 515568 328294
rect 515248 328170 515318 328226
rect 515374 328170 515442 328226
rect 515498 328170 515568 328226
rect 515248 328102 515568 328170
rect 515248 328046 515318 328102
rect 515374 328046 515442 328102
rect 515498 328046 515568 328102
rect 515248 327978 515568 328046
rect 515248 327922 515318 327978
rect 515374 327922 515442 327978
rect 515498 327922 515568 327978
rect 515248 327888 515568 327922
rect 545968 328350 546288 328384
rect 545968 328294 546038 328350
rect 546094 328294 546162 328350
rect 546218 328294 546288 328350
rect 545968 328226 546288 328294
rect 545968 328170 546038 328226
rect 546094 328170 546162 328226
rect 546218 328170 546288 328226
rect 545968 328102 546288 328170
rect 545968 328046 546038 328102
rect 546094 328046 546162 328102
rect 546218 328046 546288 328102
rect 545968 327978 546288 328046
rect 545968 327922 546038 327978
rect 546094 327922 546162 327978
rect 546218 327922 546288 327978
rect 545968 327888 546288 327922
rect 561154 328350 561774 345922
rect 561154 328294 561250 328350
rect 561306 328294 561374 328350
rect 561430 328294 561498 328350
rect 561554 328294 561622 328350
rect 561678 328294 561774 328350
rect 561154 328226 561774 328294
rect 561154 328170 561250 328226
rect 561306 328170 561374 328226
rect 561430 328170 561498 328226
rect 561554 328170 561622 328226
rect 561678 328170 561774 328226
rect 561154 328102 561774 328170
rect 561154 328046 561250 328102
rect 561306 328046 561374 328102
rect 561430 328046 561498 328102
rect 561554 328046 561622 328102
rect 561678 328046 561774 328102
rect 561154 327978 561774 328046
rect 561154 327922 561250 327978
rect 561306 327922 561374 327978
rect 561430 327922 561498 327978
rect 561554 327922 561622 327978
rect 561678 327922 561774 327978
rect 131248 316350 131568 316384
rect 131248 316294 131318 316350
rect 131374 316294 131442 316350
rect 131498 316294 131568 316350
rect 131248 316226 131568 316294
rect 131248 316170 131318 316226
rect 131374 316170 131442 316226
rect 131498 316170 131568 316226
rect 131248 316102 131568 316170
rect 131248 316046 131318 316102
rect 131374 316046 131442 316102
rect 131498 316046 131568 316102
rect 131248 315978 131568 316046
rect 131248 315922 131318 315978
rect 131374 315922 131442 315978
rect 131498 315922 131568 315978
rect 131248 315888 131568 315922
rect 161968 316350 162288 316384
rect 161968 316294 162038 316350
rect 162094 316294 162162 316350
rect 162218 316294 162288 316350
rect 161968 316226 162288 316294
rect 161968 316170 162038 316226
rect 162094 316170 162162 316226
rect 162218 316170 162288 316226
rect 161968 316102 162288 316170
rect 161968 316046 162038 316102
rect 162094 316046 162162 316102
rect 162218 316046 162288 316102
rect 161968 315978 162288 316046
rect 161968 315922 162038 315978
rect 162094 315922 162162 315978
rect 162218 315922 162288 315978
rect 161968 315888 162288 315922
rect 192688 316350 193008 316384
rect 192688 316294 192758 316350
rect 192814 316294 192882 316350
rect 192938 316294 193008 316350
rect 192688 316226 193008 316294
rect 192688 316170 192758 316226
rect 192814 316170 192882 316226
rect 192938 316170 193008 316226
rect 192688 316102 193008 316170
rect 192688 316046 192758 316102
rect 192814 316046 192882 316102
rect 192938 316046 193008 316102
rect 192688 315978 193008 316046
rect 192688 315922 192758 315978
rect 192814 315922 192882 315978
rect 192938 315922 193008 315978
rect 192688 315888 193008 315922
rect 223408 316350 223728 316384
rect 223408 316294 223478 316350
rect 223534 316294 223602 316350
rect 223658 316294 223728 316350
rect 223408 316226 223728 316294
rect 223408 316170 223478 316226
rect 223534 316170 223602 316226
rect 223658 316170 223728 316226
rect 223408 316102 223728 316170
rect 223408 316046 223478 316102
rect 223534 316046 223602 316102
rect 223658 316046 223728 316102
rect 223408 315978 223728 316046
rect 223408 315922 223478 315978
rect 223534 315922 223602 315978
rect 223658 315922 223728 315978
rect 223408 315888 223728 315922
rect 254128 316350 254448 316384
rect 254128 316294 254198 316350
rect 254254 316294 254322 316350
rect 254378 316294 254448 316350
rect 254128 316226 254448 316294
rect 254128 316170 254198 316226
rect 254254 316170 254322 316226
rect 254378 316170 254448 316226
rect 254128 316102 254448 316170
rect 254128 316046 254198 316102
rect 254254 316046 254322 316102
rect 254378 316046 254448 316102
rect 254128 315978 254448 316046
rect 254128 315922 254198 315978
rect 254254 315922 254322 315978
rect 254378 315922 254448 315978
rect 254128 315888 254448 315922
rect 284848 316350 285168 316384
rect 284848 316294 284918 316350
rect 284974 316294 285042 316350
rect 285098 316294 285168 316350
rect 284848 316226 285168 316294
rect 284848 316170 284918 316226
rect 284974 316170 285042 316226
rect 285098 316170 285168 316226
rect 284848 316102 285168 316170
rect 284848 316046 284918 316102
rect 284974 316046 285042 316102
rect 285098 316046 285168 316102
rect 284848 315978 285168 316046
rect 284848 315922 284918 315978
rect 284974 315922 285042 315978
rect 285098 315922 285168 315978
rect 284848 315888 285168 315922
rect 315568 316350 315888 316384
rect 315568 316294 315638 316350
rect 315694 316294 315762 316350
rect 315818 316294 315888 316350
rect 315568 316226 315888 316294
rect 315568 316170 315638 316226
rect 315694 316170 315762 316226
rect 315818 316170 315888 316226
rect 315568 316102 315888 316170
rect 315568 316046 315638 316102
rect 315694 316046 315762 316102
rect 315818 316046 315888 316102
rect 315568 315978 315888 316046
rect 315568 315922 315638 315978
rect 315694 315922 315762 315978
rect 315818 315922 315888 315978
rect 315568 315888 315888 315922
rect 346288 316350 346608 316384
rect 346288 316294 346358 316350
rect 346414 316294 346482 316350
rect 346538 316294 346608 316350
rect 346288 316226 346608 316294
rect 346288 316170 346358 316226
rect 346414 316170 346482 316226
rect 346538 316170 346608 316226
rect 346288 316102 346608 316170
rect 346288 316046 346358 316102
rect 346414 316046 346482 316102
rect 346538 316046 346608 316102
rect 346288 315978 346608 316046
rect 346288 315922 346358 315978
rect 346414 315922 346482 315978
rect 346538 315922 346608 315978
rect 346288 315888 346608 315922
rect 377008 316350 377328 316384
rect 377008 316294 377078 316350
rect 377134 316294 377202 316350
rect 377258 316294 377328 316350
rect 377008 316226 377328 316294
rect 377008 316170 377078 316226
rect 377134 316170 377202 316226
rect 377258 316170 377328 316226
rect 377008 316102 377328 316170
rect 377008 316046 377078 316102
rect 377134 316046 377202 316102
rect 377258 316046 377328 316102
rect 377008 315978 377328 316046
rect 377008 315922 377078 315978
rect 377134 315922 377202 315978
rect 377258 315922 377328 315978
rect 377008 315888 377328 315922
rect 407728 316350 408048 316384
rect 407728 316294 407798 316350
rect 407854 316294 407922 316350
rect 407978 316294 408048 316350
rect 407728 316226 408048 316294
rect 407728 316170 407798 316226
rect 407854 316170 407922 316226
rect 407978 316170 408048 316226
rect 407728 316102 408048 316170
rect 407728 316046 407798 316102
rect 407854 316046 407922 316102
rect 407978 316046 408048 316102
rect 407728 315978 408048 316046
rect 407728 315922 407798 315978
rect 407854 315922 407922 315978
rect 407978 315922 408048 315978
rect 407728 315888 408048 315922
rect 438448 316350 438768 316384
rect 438448 316294 438518 316350
rect 438574 316294 438642 316350
rect 438698 316294 438768 316350
rect 438448 316226 438768 316294
rect 438448 316170 438518 316226
rect 438574 316170 438642 316226
rect 438698 316170 438768 316226
rect 438448 316102 438768 316170
rect 438448 316046 438518 316102
rect 438574 316046 438642 316102
rect 438698 316046 438768 316102
rect 438448 315978 438768 316046
rect 438448 315922 438518 315978
rect 438574 315922 438642 315978
rect 438698 315922 438768 315978
rect 438448 315888 438768 315922
rect 469168 316350 469488 316384
rect 469168 316294 469238 316350
rect 469294 316294 469362 316350
rect 469418 316294 469488 316350
rect 469168 316226 469488 316294
rect 469168 316170 469238 316226
rect 469294 316170 469362 316226
rect 469418 316170 469488 316226
rect 469168 316102 469488 316170
rect 469168 316046 469238 316102
rect 469294 316046 469362 316102
rect 469418 316046 469488 316102
rect 469168 315978 469488 316046
rect 469168 315922 469238 315978
rect 469294 315922 469362 315978
rect 469418 315922 469488 315978
rect 469168 315888 469488 315922
rect 499888 316350 500208 316384
rect 499888 316294 499958 316350
rect 500014 316294 500082 316350
rect 500138 316294 500208 316350
rect 499888 316226 500208 316294
rect 499888 316170 499958 316226
rect 500014 316170 500082 316226
rect 500138 316170 500208 316226
rect 499888 316102 500208 316170
rect 499888 316046 499958 316102
rect 500014 316046 500082 316102
rect 500138 316046 500208 316102
rect 499888 315978 500208 316046
rect 499888 315922 499958 315978
rect 500014 315922 500082 315978
rect 500138 315922 500208 315978
rect 499888 315888 500208 315922
rect 530608 316350 530928 316384
rect 530608 316294 530678 316350
rect 530734 316294 530802 316350
rect 530858 316294 530928 316350
rect 530608 316226 530928 316294
rect 530608 316170 530678 316226
rect 530734 316170 530802 316226
rect 530858 316170 530928 316226
rect 530608 316102 530928 316170
rect 530608 316046 530678 316102
rect 530734 316046 530802 316102
rect 530858 316046 530928 316102
rect 530608 315978 530928 316046
rect 530608 315922 530678 315978
rect 530734 315922 530802 315978
rect 530858 315922 530928 315978
rect 530608 315888 530928 315922
rect 111154 310294 111250 310350
rect 111306 310294 111374 310350
rect 111430 310294 111498 310350
rect 111554 310294 111622 310350
rect 111678 310294 111774 310350
rect 111154 310226 111774 310294
rect 111154 310170 111250 310226
rect 111306 310170 111374 310226
rect 111430 310170 111498 310226
rect 111554 310170 111622 310226
rect 111678 310170 111774 310226
rect 111154 310102 111774 310170
rect 111154 310046 111250 310102
rect 111306 310046 111374 310102
rect 111430 310046 111498 310102
rect 111554 310046 111622 310102
rect 111678 310046 111774 310102
rect 111154 309978 111774 310046
rect 111154 309922 111250 309978
rect 111306 309922 111374 309978
rect 111430 309922 111498 309978
rect 111554 309922 111622 309978
rect 111678 309922 111774 309978
rect 96874 298294 96970 298350
rect 97026 298294 97094 298350
rect 97150 298294 97218 298350
rect 97274 298294 97342 298350
rect 97398 298294 97494 298350
rect 96874 298226 97494 298294
rect 96874 298170 96970 298226
rect 97026 298170 97094 298226
rect 97150 298170 97218 298226
rect 97274 298170 97342 298226
rect 97398 298170 97494 298226
rect 96874 298102 97494 298170
rect 96874 298046 96970 298102
rect 97026 298046 97094 298102
rect 97150 298046 97218 298102
rect 97274 298046 97342 298102
rect 97398 298046 97494 298102
rect 96874 297978 97494 298046
rect 96874 297922 96970 297978
rect 97026 297922 97094 297978
rect 97150 297922 97218 297978
rect 97274 297922 97342 297978
rect 97398 297922 97494 297978
rect 96874 280350 97494 297922
rect 100528 298350 100848 298384
rect 100528 298294 100598 298350
rect 100654 298294 100722 298350
rect 100778 298294 100848 298350
rect 100528 298226 100848 298294
rect 100528 298170 100598 298226
rect 100654 298170 100722 298226
rect 100778 298170 100848 298226
rect 100528 298102 100848 298170
rect 100528 298046 100598 298102
rect 100654 298046 100722 298102
rect 100778 298046 100848 298102
rect 100528 297978 100848 298046
rect 100528 297922 100598 297978
rect 100654 297922 100722 297978
rect 100778 297922 100848 297978
rect 100528 297888 100848 297922
rect 111154 292350 111774 309922
rect 115888 310350 116208 310384
rect 115888 310294 115958 310350
rect 116014 310294 116082 310350
rect 116138 310294 116208 310350
rect 115888 310226 116208 310294
rect 115888 310170 115958 310226
rect 116014 310170 116082 310226
rect 116138 310170 116208 310226
rect 115888 310102 116208 310170
rect 115888 310046 115958 310102
rect 116014 310046 116082 310102
rect 116138 310046 116208 310102
rect 115888 309978 116208 310046
rect 115888 309922 115958 309978
rect 116014 309922 116082 309978
rect 116138 309922 116208 309978
rect 115888 309888 116208 309922
rect 146608 310350 146928 310384
rect 146608 310294 146678 310350
rect 146734 310294 146802 310350
rect 146858 310294 146928 310350
rect 146608 310226 146928 310294
rect 146608 310170 146678 310226
rect 146734 310170 146802 310226
rect 146858 310170 146928 310226
rect 146608 310102 146928 310170
rect 146608 310046 146678 310102
rect 146734 310046 146802 310102
rect 146858 310046 146928 310102
rect 146608 309978 146928 310046
rect 146608 309922 146678 309978
rect 146734 309922 146802 309978
rect 146858 309922 146928 309978
rect 146608 309888 146928 309922
rect 177328 310350 177648 310384
rect 177328 310294 177398 310350
rect 177454 310294 177522 310350
rect 177578 310294 177648 310350
rect 177328 310226 177648 310294
rect 177328 310170 177398 310226
rect 177454 310170 177522 310226
rect 177578 310170 177648 310226
rect 177328 310102 177648 310170
rect 177328 310046 177398 310102
rect 177454 310046 177522 310102
rect 177578 310046 177648 310102
rect 177328 309978 177648 310046
rect 177328 309922 177398 309978
rect 177454 309922 177522 309978
rect 177578 309922 177648 309978
rect 177328 309888 177648 309922
rect 208048 310350 208368 310384
rect 208048 310294 208118 310350
rect 208174 310294 208242 310350
rect 208298 310294 208368 310350
rect 208048 310226 208368 310294
rect 208048 310170 208118 310226
rect 208174 310170 208242 310226
rect 208298 310170 208368 310226
rect 208048 310102 208368 310170
rect 208048 310046 208118 310102
rect 208174 310046 208242 310102
rect 208298 310046 208368 310102
rect 208048 309978 208368 310046
rect 208048 309922 208118 309978
rect 208174 309922 208242 309978
rect 208298 309922 208368 309978
rect 208048 309888 208368 309922
rect 238768 310350 239088 310384
rect 238768 310294 238838 310350
rect 238894 310294 238962 310350
rect 239018 310294 239088 310350
rect 238768 310226 239088 310294
rect 238768 310170 238838 310226
rect 238894 310170 238962 310226
rect 239018 310170 239088 310226
rect 238768 310102 239088 310170
rect 238768 310046 238838 310102
rect 238894 310046 238962 310102
rect 239018 310046 239088 310102
rect 238768 309978 239088 310046
rect 238768 309922 238838 309978
rect 238894 309922 238962 309978
rect 239018 309922 239088 309978
rect 238768 309888 239088 309922
rect 269488 310350 269808 310384
rect 269488 310294 269558 310350
rect 269614 310294 269682 310350
rect 269738 310294 269808 310350
rect 269488 310226 269808 310294
rect 269488 310170 269558 310226
rect 269614 310170 269682 310226
rect 269738 310170 269808 310226
rect 269488 310102 269808 310170
rect 269488 310046 269558 310102
rect 269614 310046 269682 310102
rect 269738 310046 269808 310102
rect 269488 309978 269808 310046
rect 269488 309922 269558 309978
rect 269614 309922 269682 309978
rect 269738 309922 269808 309978
rect 269488 309888 269808 309922
rect 300208 310350 300528 310384
rect 300208 310294 300278 310350
rect 300334 310294 300402 310350
rect 300458 310294 300528 310350
rect 300208 310226 300528 310294
rect 300208 310170 300278 310226
rect 300334 310170 300402 310226
rect 300458 310170 300528 310226
rect 300208 310102 300528 310170
rect 300208 310046 300278 310102
rect 300334 310046 300402 310102
rect 300458 310046 300528 310102
rect 300208 309978 300528 310046
rect 300208 309922 300278 309978
rect 300334 309922 300402 309978
rect 300458 309922 300528 309978
rect 300208 309888 300528 309922
rect 330928 310350 331248 310384
rect 330928 310294 330998 310350
rect 331054 310294 331122 310350
rect 331178 310294 331248 310350
rect 330928 310226 331248 310294
rect 330928 310170 330998 310226
rect 331054 310170 331122 310226
rect 331178 310170 331248 310226
rect 330928 310102 331248 310170
rect 330928 310046 330998 310102
rect 331054 310046 331122 310102
rect 331178 310046 331248 310102
rect 330928 309978 331248 310046
rect 330928 309922 330998 309978
rect 331054 309922 331122 309978
rect 331178 309922 331248 309978
rect 330928 309888 331248 309922
rect 361648 310350 361968 310384
rect 361648 310294 361718 310350
rect 361774 310294 361842 310350
rect 361898 310294 361968 310350
rect 361648 310226 361968 310294
rect 361648 310170 361718 310226
rect 361774 310170 361842 310226
rect 361898 310170 361968 310226
rect 361648 310102 361968 310170
rect 361648 310046 361718 310102
rect 361774 310046 361842 310102
rect 361898 310046 361968 310102
rect 361648 309978 361968 310046
rect 361648 309922 361718 309978
rect 361774 309922 361842 309978
rect 361898 309922 361968 309978
rect 361648 309888 361968 309922
rect 392368 310350 392688 310384
rect 392368 310294 392438 310350
rect 392494 310294 392562 310350
rect 392618 310294 392688 310350
rect 392368 310226 392688 310294
rect 392368 310170 392438 310226
rect 392494 310170 392562 310226
rect 392618 310170 392688 310226
rect 392368 310102 392688 310170
rect 392368 310046 392438 310102
rect 392494 310046 392562 310102
rect 392618 310046 392688 310102
rect 392368 309978 392688 310046
rect 392368 309922 392438 309978
rect 392494 309922 392562 309978
rect 392618 309922 392688 309978
rect 392368 309888 392688 309922
rect 423088 310350 423408 310384
rect 423088 310294 423158 310350
rect 423214 310294 423282 310350
rect 423338 310294 423408 310350
rect 423088 310226 423408 310294
rect 423088 310170 423158 310226
rect 423214 310170 423282 310226
rect 423338 310170 423408 310226
rect 423088 310102 423408 310170
rect 423088 310046 423158 310102
rect 423214 310046 423282 310102
rect 423338 310046 423408 310102
rect 423088 309978 423408 310046
rect 423088 309922 423158 309978
rect 423214 309922 423282 309978
rect 423338 309922 423408 309978
rect 423088 309888 423408 309922
rect 453808 310350 454128 310384
rect 453808 310294 453878 310350
rect 453934 310294 454002 310350
rect 454058 310294 454128 310350
rect 453808 310226 454128 310294
rect 453808 310170 453878 310226
rect 453934 310170 454002 310226
rect 454058 310170 454128 310226
rect 453808 310102 454128 310170
rect 453808 310046 453878 310102
rect 453934 310046 454002 310102
rect 454058 310046 454128 310102
rect 453808 309978 454128 310046
rect 453808 309922 453878 309978
rect 453934 309922 454002 309978
rect 454058 309922 454128 309978
rect 453808 309888 454128 309922
rect 484528 310350 484848 310384
rect 484528 310294 484598 310350
rect 484654 310294 484722 310350
rect 484778 310294 484848 310350
rect 484528 310226 484848 310294
rect 484528 310170 484598 310226
rect 484654 310170 484722 310226
rect 484778 310170 484848 310226
rect 484528 310102 484848 310170
rect 484528 310046 484598 310102
rect 484654 310046 484722 310102
rect 484778 310046 484848 310102
rect 484528 309978 484848 310046
rect 484528 309922 484598 309978
rect 484654 309922 484722 309978
rect 484778 309922 484848 309978
rect 484528 309888 484848 309922
rect 515248 310350 515568 310384
rect 515248 310294 515318 310350
rect 515374 310294 515442 310350
rect 515498 310294 515568 310350
rect 515248 310226 515568 310294
rect 515248 310170 515318 310226
rect 515374 310170 515442 310226
rect 515498 310170 515568 310226
rect 515248 310102 515568 310170
rect 515248 310046 515318 310102
rect 515374 310046 515442 310102
rect 515498 310046 515568 310102
rect 515248 309978 515568 310046
rect 515248 309922 515318 309978
rect 515374 309922 515442 309978
rect 515498 309922 515568 309978
rect 515248 309888 515568 309922
rect 545968 310350 546288 310384
rect 545968 310294 546038 310350
rect 546094 310294 546162 310350
rect 546218 310294 546288 310350
rect 545968 310226 546288 310294
rect 545968 310170 546038 310226
rect 546094 310170 546162 310226
rect 546218 310170 546288 310226
rect 545968 310102 546288 310170
rect 545968 310046 546038 310102
rect 546094 310046 546162 310102
rect 546218 310046 546288 310102
rect 545968 309978 546288 310046
rect 545968 309922 546038 309978
rect 546094 309922 546162 309978
rect 546218 309922 546288 309978
rect 545968 309888 546288 309922
rect 561154 310350 561774 327922
rect 561154 310294 561250 310350
rect 561306 310294 561374 310350
rect 561430 310294 561498 310350
rect 561554 310294 561622 310350
rect 561678 310294 561774 310350
rect 561154 310226 561774 310294
rect 561154 310170 561250 310226
rect 561306 310170 561374 310226
rect 561430 310170 561498 310226
rect 561554 310170 561622 310226
rect 561678 310170 561774 310226
rect 561154 310102 561774 310170
rect 561154 310046 561250 310102
rect 561306 310046 561374 310102
rect 561430 310046 561498 310102
rect 561554 310046 561622 310102
rect 561678 310046 561774 310102
rect 561154 309978 561774 310046
rect 561154 309922 561250 309978
rect 561306 309922 561374 309978
rect 561430 309922 561498 309978
rect 561554 309922 561622 309978
rect 561678 309922 561774 309978
rect 131248 298350 131568 298384
rect 131248 298294 131318 298350
rect 131374 298294 131442 298350
rect 131498 298294 131568 298350
rect 131248 298226 131568 298294
rect 131248 298170 131318 298226
rect 131374 298170 131442 298226
rect 131498 298170 131568 298226
rect 131248 298102 131568 298170
rect 131248 298046 131318 298102
rect 131374 298046 131442 298102
rect 131498 298046 131568 298102
rect 131248 297978 131568 298046
rect 131248 297922 131318 297978
rect 131374 297922 131442 297978
rect 131498 297922 131568 297978
rect 131248 297888 131568 297922
rect 161968 298350 162288 298384
rect 161968 298294 162038 298350
rect 162094 298294 162162 298350
rect 162218 298294 162288 298350
rect 161968 298226 162288 298294
rect 161968 298170 162038 298226
rect 162094 298170 162162 298226
rect 162218 298170 162288 298226
rect 161968 298102 162288 298170
rect 161968 298046 162038 298102
rect 162094 298046 162162 298102
rect 162218 298046 162288 298102
rect 161968 297978 162288 298046
rect 161968 297922 162038 297978
rect 162094 297922 162162 297978
rect 162218 297922 162288 297978
rect 161968 297888 162288 297922
rect 192688 298350 193008 298384
rect 192688 298294 192758 298350
rect 192814 298294 192882 298350
rect 192938 298294 193008 298350
rect 192688 298226 193008 298294
rect 192688 298170 192758 298226
rect 192814 298170 192882 298226
rect 192938 298170 193008 298226
rect 192688 298102 193008 298170
rect 192688 298046 192758 298102
rect 192814 298046 192882 298102
rect 192938 298046 193008 298102
rect 192688 297978 193008 298046
rect 192688 297922 192758 297978
rect 192814 297922 192882 297978
rect 192938 297922 193008 297978
rect 192688 297888 193008 297922
rect 223408 298350 223728 298384
rect 223408 298294 223478 298350
rect 223534 298294 223602 298350
rect 223658 298294 223728 298350
rect 223408 298226 223728 298294
rect 223408 298170 223478 298226
rect 223534 298170 223602 298226
rect 223658 298170 223728 298226
rect 223408 298102 223728 298170
rect 223408 298046 223478 298102
rect 223534 298046 223602 298102
rect 223658 298046 223728 298102
rect 223408 297978 223728 298046
rect 223408 297922 223478 297978
rect 223534 297922 223602 297978
rect 223658 297922 223728 297978
rect 223408 297888 223728 297922
rect 254128 298350 254448 298384
rect 254128 298294 254198 298350
rect 254254 298294 254322 298350
rect 254378 298294 254448 298350
rect 254128 298226 254448 298294
rect 254128 298170 254198 298226
rect 254254 298170 254322 298226
rect 254378 298170 254448 298226
rect 254128 298102 254448 298170
rect 254128 298046 254198 298102
rect 254254 298046 254322 298102
rect 254378 298046 254448 298102
rect 254128 297978 254448 298046
rect 254128 297922 254198 297978
rect 254254 297922 254322 297978
rect 254378 297922 254448 297978
rect 254128 297888 254448 297922
rect 284848 298350 285168 298384
rect 284848 298294 284918 298350
rect 284974 298294 285042 298350
rect 285098 298294 285168 298350
rect 284848 298226 285168 298294
rect 284848 298170 284918 298226
rect 284974 298170 285042 298226
rect 285098 298170 285168 298226
rect 284848 298102 285168 298170
rect 284848 298046 284918 298102
rect 284974 298046 285042 298102
rect 285098 298046 285168 298102
rect 284848 297978 285168 298046
rect 284848 297922 284918 297978
rect 284974 297922 285042 297978
rect 285098 297922 285168 297978
rect 284848 297888 285168 297922
rect 315568 298350 315888 298384
rect 315568 298294 315638 298350
rect 315694 298294 315762 298350
rect 315818 298294 315888 298350
rect 315568 298226 315888 298294
rect 315568 298170 315638 298226
rect 315694 298170 315762 298226
rect 315818 298170 315888 298226
rect 315568 298102 315888 298170
rect 315568 298046 315638 298102
rect 315694 298046 315762 298102
rect 315818 298046 315888 298102
rect 315568 297978 315888 298046
rect 315568 297922 315638 297978
rect 315694 297922 315762 297978
rect 315818 297922 315888 297978
rect 315568 297888 315888 297922
rect 346288 298350 346608 298384
rect 346288 298294 346358 298350
rect 346414 298294 346482 298350
rect 346538 298294 346608 298350
rect 346288 298226 346608 298294
rect 346288 298170 346358 298226
rect 346414 298170 346482 298226
rect 346538 298170 346608 298226
rect 346288 298102 346608 298170
rect 346288 298046 346358 298102
rect 346414 298046 346482 298102
rect 346538 298046 346608 298102
rect 346288 297978 346608 298046
rect 346288 297922 346358 297978
rect 346414 297922 346482 297978
rect 346538 297922 346608 297978
rect 346288 297888 346608 297922
rect 377008 298350 377328 298384
rect 377008 298294 377078 298350
rect 377134 298294 377202 298350
rect 377258 298294 377328 298350
rect 377008 298226 377328 298294
rect 377008 298170 377078 298226
rect 377134 298170 377202 298226
rect 377258 298170 377328 298226
rect 377008 298102 377328 298170
rect 377008 298046 377078 298102
rect 377134 298046 377202 298102
rect 377258 298046 377328 298102
rect 377008 297978 377328 298046
rect 377008 297922 377078 297978
rect 377134 297922 377202 297978
rect 377258 297922 377328 297978
rect 377008 297888 377328 297922
rect 407728 298350 408048 298384
rect 407728 298294 407798 298350
rect 407854 298294 407922 298350
rect 407978 298294 408048 298350
rect 407728 298226 408048 298294
rect 407728 298170 407798 298226
rect 407854 298170 407922 298226
rect 407978 298170 408048 298226
rect 407728 298102 408048 298170
rect 407728 298046 407798 298102
rect 407854 298046 407922 298102
rect 407978 298046 408048 298102
rect 407728 297978 408048 298046
rect 407728 297922 407798 297978
rect 407854 297922 407922 297978
rect 407978 297922 408048 297978
rect 407728 297888 408048 297922
rect 438448 298350 438768 298384
rect 438448 298294 438518 298350
rect 438574 298294 438642 298350
rect 438698 298294 438768 298350
rect 438448 298226 438768 298294
rect 438448 298170 438518 298226
rect 438574 298170 438642 298226
rect 438698 298170 438768 298226
rect 438448 298102 438768 298170
rect 438448 298046 438518 298102
rect 438574 298046 438642 298102
rect 438698 298046 438768 298102
rect 438448 297978 438768 298046
rect 438448 297922 438518 297978
rect 438574 297922 438642 297978
rect 438698 297922 438768 297978
rect 438448 297888 438768 297922
rect 469168 298350 469488 298384
rect 469168 298294 469238 298350
rect 469294 298294 469362 298350
rect 469418 298294 469488 298350
rect 469168 298226 469488 298294
rect 469168 298170 469238 298226
rect 469294 298170 469362 298226
rect 469418 298170 469488 298226
rect 469168 298102 469488 298170
rect 469168 298046 469238 298102
rect 469294 298046 469362 298102
rect 469418 298046 469488 298102
rect 469168 297978 469488 298046
rect 469168 297922 469238 297978
rect 469294 297922 469362 297978
rect 469418 297922 469488 297978
rect 469168 297888 469488 297922
rect 499888 298350 500208 298384
rect 499888 298294 499958 298350
rect 500014 298294 500082 298350
rect 500138 298294 500208 298350
rect 499888 298226 500208 298294
rect 499888 298170 499958 298226
rect 500014 298170 500082 298226
rect 500138 298170 500208 298226
rect 499888 298102 500208 298170
rect 499888 298046 499958 298102
rect 500014 298046 500082 298102
rect 500138 298046 500208 298102
rect 499888 297978 500208 298046
rect 499888 297922 499958 297978
rect 500014 297922 500082 297978
rect 500138 297922 500208 297978
rect 499888 297888 500208 297922
rect 530608 298350 530928 298384
rect 530608 298294 530678 298350
rect 530734 298294 530802 298350
rect 530858 298294 530928 298350
rect 530608 298226 530928 298294
rect 530608 298170 530678 298226
rect 530734 298170 530802 298226
rect 530858 298170 530928 298226
rect 530608 298102 530928 298170
rect 530608 298046 530678 298102
rect 530734 298046 530802 298102
rect 530858 298046 530928 298102
rect 530608 297978 530928 298046
rect 530608 297922 530678 297978
rect 530734 297922 530802 297978
rect 530858 297922 530928 297978
rect 530608 297888 530928 297922
rect 111154 292294 111250 292350
rect 111306 292294 111374 292350
rect 111430 292294 111498 292350
rect 111554 292294 111622 292350
rect 111678 292294 111774 292350
rect 111154 292226 111774 292294
rect 111154 292170 111250 292226
rect 111306 292170 111374 292226
rect 111430 292170 111498 292226
rect 111554 292170 111622 292226
rect 111678 292170 111774 292226
rect 111154 292102 111774 292170
rect 111154 292046 111250 292102
rect 111306 292046 111374 292102
rect 111430 292046 111498 292102
rect 111554 292046 111622 292102
rect 111678 292046 111774 292102
rect 111154 291978 111774 292046
rect 111154 291922 111250 291978
rect 111306 291922 111374 291978
rect 111430 291922 111498 291978
rect 111554 291922 111622 291978
rect 111678 291922 111774 291978
rect 96874 280294 96970 280350
rect 97026 280294 97094 280350
rect 97150 280294 97218 280350
rect 97274 280294 97342 280350
rect 97398 280294 97494 280350
rect 96874 280226 97494 280294
rect 96874 280170 96970 280226
rect 97026 280170 97094 280226
rect 97150 280170 97218 280226
rect 97274 280170 97342 280226
rect 97398 280170 97494 280226
rect 96874 280102 97494 280170
rect 96874 280046 96970 280102
rect 97026 280046 97094 280102
rect 97150 280046 97218 280102
rect 97274 280046 97342 280102
rect 97398 280046 97494 280102
rect 96874 279978 97494 280046
rect 96874 279922 96970 279978
rect 97026 279922 97094 279978
rect 97150 279922 97218 279978
rect 97274 279922 97342 279978
rect 97398 279922 97494 279978
rect 96874 262350 97494 279922
rect 100528 280350 100848 280384
rect 100528 280294 100598 280350
rect 100654 280294 100722 280350
rect 100778 280294 100848 280350
rect 100528 280226 100848 280294
rect 100528 280170 100598 280226
rect 100654 280170 100722 280226
rect 100778 280170 100848 280226
rect 100528 280102 100848 280170
rect 100528 280046 100598 280102
rect 100654 280046 100722 280102
rect 100778 280046 100848 280102
rect 100528 279978 100848 280046
rect 100528 279922 100598 279978
rect 100654 279922 100722 279978
rect 100778 279922 100848 279978
rect 100528 279888 100848 279922
rect 111154 274350 111774 291922
rect 115888 292350 116208 292384
rect 115888 292294 115958 292350
rect 116014 292294 116082 292350
rect 116138 292294 116208 292350
rect 115888 292226 116208 292294
rect 115888 292170 115958 292226
rect 116014 292170 116082 292226
rect 116138 292170 116208 292226
rect 115888 292102 116208 292170
rect 115888 292046 115958 292102
rect 116014 292046 116082 292102
rect 116138 292046 116208 292102
rect 115888 291978 116208 292046
rect 115888 291922 115958 291978
rect 116014 291922 116082 291978
rect 116138 291922 116208 291978
rect 115888 291888 116208 291922
rect 146608 292350 146928 292384
rect 146608 292294 146678 292350
rect 146734 292294 146802 292350
rect 146858 292294 146928 292350
rect 146608 292226 146928 292294
rect 146608 292170 146678 292226
rect 146734 292170 146802 292226
rect 146858 292170 146928 292226
rect 146608 292102 146928 292170
rect 146608 292046 146678 292102
rect 146734 292046 146802 292102
rect 146858 292046 146928 292102
rect 146608 291978 146928 292046
rect 146608 291922 146678 291978
rect 146734 291922 146802 291978
rect 146858 291922 146928 291978
rect 146608 291888 146928 291922
rect 177328 292350 177648 292384
rect 177328 292294 177398 292350
rect 177454 292294 177522 292350
rect 177578 292294 177648 292350
rect 177328 292226 177648 292294
rect 177328 292170 177398 292226
rect 177454 292170 177522 292226
rect 177578 292170 177648 292226
rect 177328 292102 177648 292170
rect 177328 292046 177398 292102
rect 177454 292046 177522 292102
rect 177578 292046 177648 292102
rect 177328 291978 177648 292046
rect 177328 291922 177398 291978
rect 177454 291922 177522 291978
rect 177578 291922 177648 291978
rect 177328 291888 177648 291922
rect 208048 292350 208368 292384
rect 208048 292294 208118 292350
rect 208174 292294 208242 292350
rect 208298 292294 208368 292350
rect 208048 292226 208368 292294
rect 208048 292170 208118 292226
rect 208174 292170 208242 292226
rect 208298 292170 208368 292226
rect 208048 292102 208368 292170
rect 208048 292046 208118 292102
rect 208174 292046 208242 292102
rect 208298 292046 208368 292102
rect 208048 291978 208368 292046
rect 208048 291922 208118 291978
rect 208174 291922 208242 291978
rect 208298 291922 208368 291978
rect 208048 291888 208368 291922
rect 238768 292350 239088 292384
rect 238768 292294 238838 292350
rect 238894 292294 238962 292350
rect 239018 292294 239088 292350
rect 238768 292226 239088 292294
rect 238768 292170 238838 292226
rect 238894 292170 238962 292226
rect 239018 292170 239088 292226
rect 238768 292102 239088 292170
rect 238768 292046 238838 292102
rect 238894 292046 238962 292102
rect 239018 292046 239088 292102
rect 238768 291978 239088 292046
rect 238768 291922 238838 291978
rect 238894 291922 238962 291978
rect 239018 291922 239088 291978
rect 238768 291888 239088 291922
rect 269488 292350 269808 292384
rect 269488 292294 269558 292350
rect 269614 292294 269682 292350
rect 269738 292294 269808 292350
rect 269488 292226 269808 292294
rect 269488 292170 269558 292226
rect 269614 292170 269682 292226
rect 269738 292170 269808 292226
rect 269488 292102 269808 292170
rect 269488 292046 269558 292102
rect 269614 292046 269682 292102
rect 269738 292046 269808 292102
rect 269488 291978 269808 292046
rect 269488 291922 269558 291978
rect 269614 291922 269682 291978
rect 269738 291922 269808 291978
rect 269488 291888 269808 291922
rect 300208 292350 300528 292384
rect 300208 292294 300278 292350
rect 300334 292294 300402 292350
rect 300458 292294 300528 292350
rect 300208 292226 300528 292294
rect 300208 292170 300278 292226
rect 300334 292170 300402 292226
rect 300458 292170 300528 292226
rect 300208 292102 300528 292170
rect 300208 292046 300278 292102
rect 300334 292046 300402 292102
rect 300458 292046 300528 292102
rect 300208 291978 300528 292046
rect 300208 291922 300278 291978
rect 300334 291922 300402 291978
rect 300458 291922 300528 291978
rect 300208 291888 300528 291922
rect 330928 292350 331248 292384
rect 330928 292294 330998 292350
rect 331054 292294 331122 292350
rect 331178 292294 331248 292350
rect 330928 292226 331248 292294
rect 330928 292170 330998 292226
rect 331054 292170 331122 292226
rect 331178 292170 331248 292226
rect 330928 292102 331248 292170
rect 330928 292046 330998 292102
rect 331054 292046 331122 292102
rect 331178 292046 331248 292102
rect 330928 291978 331248 292046
rect 330928 291922 330998 291978
rect 331054 291922 331122 291978
rect 331178 291922 331248 291978
rect 330928 291888 331248 291922
rect 361648 292350 361968 292384
rect 361648 292294 361718 292350
rect 361774 292294 361842 292350
rect 361898 292294 361968 292350
rect 361648 292226 361968 292294
rect 361648 292170 361718 292226
rect 361774 292170 361842 292226
rect 361898 292170 361968 292226
rect 361648 292102 361968 292170
rect 361648 292046 361718 292102
rect 361774 292046 361842 292102
rect 361898 292046 361968 292102
rect 361648 291978 361968 292046
rect 361648 291922 361718 291978
rect 361774 291922 361842 291978
rect 361898 291922 361968 291978
rect 361648 291888 361968 291922
rect 392368 292350 392688 292384
rect 392368 292294 392438 292350
rect 392494 292294 392562 292350
rect 392618 292294 392688 292350
rect 392368 292226 392688 292294
rect 392368 292170 392438 292226
rect 392494 292170 392562 292226
rect 392618 292170 392688 292226
rect 392368 292102 392688 292170
rect 392368 292046 392438 292102
rect 392494 292046 392562 292102
rect 392618 292046 392688 292102
rect 392368 291978 392688 292046
rect 392368 291922 392438 291978
rect 392494 291922 392562 291978
rect 392618 291922 392688 291978
rect 392368 291888 392688 291922
rect 423088 292350 423408 292384
rect 423088 292294 423158 292350
rect 423214 292294 423282 292350
rect 423338 292294 423408 292350
rect 423088 292226 423408 292294
rect 423088 292170 423158 292226
rect 423214 292170 423282 292226
rect 423338 292170 423408 292226
rect 423088 292102 423408 292170
rect 423088 292046 423158 292102
rect 423214 292046 423282 292102
rect 423338 292046 423408 292102
rect 423088 291978 423408 292046
rect 423088 291922 423158 291978
rect 423214 291922 423282 291978
rect 423338 291922 423408 291978
rect 423088 291888 423408 291922
rect 453808 292350 454128 292384
rect 453808 292294 453878 292350
rect 453934 292294 454002 292350
rect 454058 292294 454128 292350
rect 453808 292226 454128 292294
rect 453808 292170 453878 292226
rect 453934 292170 454002 292226
rect 454058 292170 454128 292226
rect 453808 292102 454128 292170
rect 453808 292046 453878 292102
rect 453934 292046 454002 292102
rect 454058 292046 454128 292102
rect 453808 291978 454128 292046
rect 453808 291922 453878 291978
rect 453934 291922 454002 291978
rect 454058 291922 454128 291978
rect 453808 291888 454128 291922
rect 484528 292350 484848 292384
rect 484528 292294 484598 292350
rect 484654 292294 484722 292350
rect 484778 292294 484848 292350
rect 484528 292226 484848 292294
rect 484528 292170 484598 292226
rect 484654 292170 484722 292226
rect 484778 292170 484848 292226
rect 484528 292102 484848 292170
rect 484528 292046 484598 292102
rect 484654 292046 484722 292102
rect 484778 292046 484848 292102
rect 484528 291978 484848 292046
rect 484528 291922 484598 291978
rect 484654 291922 484722 291978
rect 484778 291922 484848 291978
rect 484528 291888 484848 291922
rect 515248 292350 515568 292384
rect 515248 292294 515318 292350
rect 515374 292294 515442 292350
rect 515498 292294 515568 292350
rect 515248 292226 515568 292294
rect 515248 292170 515318 292226
rect 515374 292170 515442 292226
rect 515498 292170 515568 292226
rect 515248 292102 515568 292170
rect 515248 292046 515318 292102
rect 515374 292046 515442 292102
rect 515498 292046 515568 292102
rect 515248 291978 515568 292046
rect 515248 291922 515318 291978
rect 515374 291922 515442 291978
rect 515498 291922 515568 291978
rect 515248 291888 515568 291922
rect 545968 292350 546288 292384
rect 545968 292294 546038 292350
rect 546094 292294 546162 292350
rect 546218 292294 546288 292350
rect 545968 292226 546288 292294
rect 545968 292170 546038 292226
rect 546094 292170 546162 292226
rect 546218 292170 546288 292226
rect 545968 292102 546288 292170
rect 545968 292046 546038 292102
rect 546094 292046 546162 292102
rect 546218 292046 546288 292102
rect 545968 291978 546288 292046
rect 545968 291922 546038 291978
rect 546094 291922 546162 291978
rect 546218 291922 546288 291978
rect 545968 291888 546288 291922
rect 561154 292350 561774 309922
rect 561154 292294 561250 292350
rect 561306 292294 561374 292350
rect 561430 292294 561498 292350
rect 561554 292294 561622 292350
rect 561678 292294 561774 292350
rect 561154 292226 561774 292294
rect 561154 292170 561250 292226
rect 561306 292170 561374 292226
rect 561430 292170 561498 292226
rect 561554 292170 561622 292226
rect 561678 292170 561774 292226
rect 561154 292102 561774 292170
rect 561154 292046 561250 292102
rect 561306 292046 561374 292102
rect 561430 292046 561498 292102
rect 561554 292046 561622 292102
rect 561678 292046 561774 292102
rect 561154 291978 561774 292046
rect 561154 291922 561250 291978
rect 561306 291922 561374 291978
rect 561430 291922 561498 291978
rect 561554 291922 561622 291978
rect 561678 291922 561774 291978
rect 131248 280350 131568 280384
rect 131248 280294 131318 280350
rect 131374 280294 131442 280350
rect 131498 280294 131568 280350
rect 131248 280226 131568 280294
rect 131248 280170 131318 280226
rect 131374 280170 131442 280226
rect 131498 280170 131568 280226
rect 131248 280102 131568 280170
rect 131248 280046 131318 280102
rect 131374 280046 131442 280102
rect 131498 280046 131568 280102
rect 131248 279978 131568 280046
rect 131248 279922 131318 279978
rect 131374 279922 131442 279978
rect 131498 279922 131568 279978
rect 131248 279888 131568 279922
rect 161968 280350 162288 280384
rect 161968 280294 162038 280350
rect 162094 280294 162162 280350
rect 162218 280294 162288 280350
rect 161968 280226 162288 280294
rect 161968 280170 162038 280226
rect 162094 280170 162162 280226
rect 162218 280170 162288 280226
rect 161968 280102 162288 280170
rect 161968 280046 162038 280102
rect 162094 280046 162162 280102
rect 162218 280046 162288 280102
rect 161968 279978 162288 280046
rect 161968 279922 162038 279978
rect 162094 279922 162162 279978
rect 162218 279922 162288 279978
rect 161968 279888 162288 279922
rect 192688 280350 193008 280384
rect 192688 280294 192758 280350
rect 192814 280294 192882 280350
rect 192938 280294 193008 280350
rect 192688 280226 193008 280294
rect 192688 280170 192758 280226
rect 192814 280170 192882 280226
rect 192938 280170 193008 280226
rect 192688 280102 193008 280170
rect 192688 280046 192758 280102
rect 192814 280046 192882 280102
rect 192938 280046 193008 280102
rect 192688 279978 193008 280046
rect 192688 279922 192758 279978
rect 192814 279922 192882 279978
rect 192938 279922 193008 279978
rect 192688 279888 193008 279922
rect 223408 280350 223728 280384
rect 223408 280294 223478 280350
rect 223534 280294 223602 280350
rect 223658 280294 223728 280350
rect 223408 280226 223728 280294
rect 223408 280170 223478 280226
rect 223534 280170 223602 280226
rect 223658 280170 223728 280226
rect 223408 280102 223728 280170
rect 223408 280046 223478 280102
rect 223534 280046 223602 280102
rect 223658 280046 223728 280102
rect 223408 279978 223728 280046
rect 223408 279922 223478 279978
rect 223534 279922 223602 279978
rect 223658 279922 223728 279978
rect 223408 279888 223728 279922
rect 254128 280350 254448 280384
rect 254128 280294 254198 280350
rect 254254 280294 254322 280350
rect 254378 280294 254448 280350
rect 254128 280226 254448 280294
rect 254128 280170 254198 280226
rect 254254 280170 254322 280226
rect 254378 280170 254448 280226
rect 254128 280102 254448 280170
rect 254128 280046 254198 280102
rect 254254 280046 254322 280102
rect 254378 280046 254448 280102
rect 254128 279978 254448 280046
rect 254128 279922 254198 279978
rect 254254 279922 254322 279978
rect 254378 279922 254448 279978
rect 254128 279888 254448 279922
rect 284848 280350 285168 280384
rect 284848 280294 284918 280350
rect 284974 280294 285042 280350
rect 285098 280294 285168 280350
rect 284848 280226 285168 280294
rect 284848 280170 284918 280226
rect 284974 280170 285042 280226
rect 285098 280170 285168 280226
rect 284848 280102 285168 280170
rect 284848 280046 284918 280102
rect 284974 280046 285042 280102
rect 285098 280046 285168 280102
rect 284848 279978 285168 280046
rect 284848 279922 284918 279978
rect 284974 279922 285042 279978
rect 285098 279922 285168 279978
rect 284848 279888 285168 279922
rect 315568 280350 315888 280384
rect 315568 280294 315638 280350
rect 315694 280294 315762 280350
rect 315818 280294 315888 280350
rect 315568 280226 315888 280294
rect 315568 280170 315638 280226
rect 315694 280170 315762 280226
rect 315818 280170 315888 280226
rect 315568 280102 315888 280170
rect 315568 280046 315638 280102
rect 315694 280046 315762 280102
rect 315818 280046 315888 280102
rect 315568 279978 315888 280046
rect 315568 279922 315638 279978
rect 315694 279922 315762 279978
rect 315818 279922 315888 279978
rect 315568 279888 315888 279922
rect 346288 280350 346608 280384
rect 346288 280294 346358 280350
rect 346414 280294 346482 280350
rect 346538 280294 346608 280350
rect 346288 280226 346608 280294
rect 346288 280170 346358 280226
rect 346414 280170 346482 280226
rect 346538 280170 346608 280226
rect 346288 280102 346608 280170
rect 346288 280046 346358 280102
rect 346414 280046 346482 280102
rect 346538 280046 346608 280102
rect 346288 279978 346608 280046
rect 346288 279922 346358 279978
rect 346414 279922 346482 279978
rect 346538 279922 346608 279978
rect 346288 279888 346608 279922
rect 377008 280350 377328 280384
rect 377008 280294 377078 280350
rect 377134 280294 377202 280350
rect 377258 280294 377328 280350
rect 377008 280226 377328 280294
rect 377008 280170 377078 280226
rect 377134 280170 377202 280226
rect 377258 280170 377328 280226
rect 377008 280102 377328 280170
rect 377008 280046 377078 280102
rect 377134 280046 377202 280102
rect 377258 280046 377328 280102
rect 377008 279978 377328 280046
rect 377008 279922 377078 279978
rect 377134 279922 377202 279978
rect 377258 279922 377328 279978
rect 377008 279888 377328 279922
rect 407728 280350 408048 280384
rect 407728 280294 407798 280350
rect 407854 280294 407922 280350
rect 407978 280294 408048 280350
rect 407728 280226 408048 280294
rect 407728 280170 407798 280226
rect 407854 280170 407922 280226
rect 407978 280170 408048 280226
rect 407728 280102 408048 280170
rect 407728 280046 407798 280102
rect 407854 280046 407922 280102
rect 407978 280046 408048 280102
rect 407728 279978 408048 280046
rect 407728 279922 407798 279978
rect 407854 279922 407922 279978
rect 407978 279922 408048 279978
rect 407728 279888 408048 279922
rect 438448 280350 438768 280384
rect 438448 280294 438518 280350
rect 438574 280294 438642 280350
rect 438698 280294 438768 280350
rect 438448 280226 438768 280294
rect 438448 280170 438518 280226
rect 438574 280170 438642 280226
rect 438698 280170 438768 280226
rect 438448 280102 438768 280170
rect 438448 280046 438518 280102
rect 438574 280046 438642 280102
rect 438698 280046 438768 280102
rect 438448 279978 438768 280046
rect 438448 279922 438518 279978
rect 438574 279922 438642 279978
rect 438698 279922 438768 279978
rect 438448 279888 438768 279922
rect 469168 280350 469488 280384
rect 469168 280294 469238 280350
rect 469294 280294 469362 280350
rect 469418 280294 469488 280350
rect 469168 280226 469488 280294
rect 469168 280170 469238 280226
rect 469294 280170 469362 280226
rect 469418 280170 469488 280226
rect 469168 280102 469488 280170
rect 469168 280046 469238 280102
rect 469294 280046 469362 280102
rect 469418 280046 469488 280102
rect 469168 279978 469488 280046
rect 469168 279922 469238 279978
rect 469294 279922 469362 279978
rect 469418 279922 469488 279978
rect 469168 279888 469488 279922
rect 499888 280350 500208 280384
rect 499888 280294 499958 280350
rect 500014 280294 500082 280350
rect 500138 280294 500208 280350
rect 499888 280226 500208 280294
rect 499888 280170 499958 280226
rect 500014 280170 500082 280226
rect 500138 280170 500208 280226
rect 499888 280102 500208 280170
rect 499888 280046 499958 280102
rect 500014 280046 500082 280102
rect 500138 280046 500208 280102
rect 499888 279978 500208 280046
rect 499888 279922 499958 279978
rect 500014 279922 500082 279978
rect 500138 279922 500208 279978
rect 499888 279888 500208 279922
rect 530608 280350 530928 280384
rect 530608 280294 530678 280350
rect 530734 280294 530802 280350
rect 530858 280294 530928 280350
rect 530608 280226 530928 280294
rect 530608 280170 530678 280226
rect 530734 280170 530802 280226
rect 530858 280170 530928 280226
rect 530608 280102 530928 280170
rect 530608 280046 530678 280102
rect 530734 280046 530802 280102
rect 530858 280046 530928 280102
rect 530608 279978 530928 280046
rect 530608 279922 530678 279978
rect 530734 279922 530802 279978
rect 530858 279922 530928 279978
rect 530608 279888 530928 279922
rect 111154 274294 111250 274350
rect 111306 274294 111374 274350
rect 111430 274294 111498 274350
rect 111554 274294 111622 274350
rect 111678 274294 111774 274350
rect 111154 274226 111774 274294
rect 111154 274170 111250 274226
rect 111306 274170 111374 274226
rect 111430 274170 111498 274226
rect 111554 274170 111622 274226
rect 111678 274170 111774 274226
rect 111154 274102 111774 274170
rect 111154 274046 111250 274102
rect 111306 274046 111374 274102
rect 111430 274046 111498 274102
rect 111554 274046 111622 274102
rect 111678 274046 111774 274102
rect 111154 273978 111774 274046
rect 111154 273922 111250 273978
rect 111306 273922 111374 273978
rect 111430 273922 111498 273978
rect 111554 273922 111622 273978
rect 111678 273922 111774 273978
rect 96874 262294 96970 262350
rect 97026 262294 97094 262350
rect 97150 262294 97218 262350
rect 97274 262294 97342 262350
rect 97398 262294 97494 262350
rect 96874 262226 97494 262294
rect 96874 262170 96970 262226
rect 97026 262170 97094 262226
rect 97150 262170 97218 262226
rect 97274 262170 97342 262226
rect 97398 262170 97494 262226
rect 96874 262102 97494 262170
rect 96874 262046 96970 262102
rect 97026 262046 97094 262102
rect 97150 262046 97218 262102
rect 97274 262046 97342 262102
rect 97398 262046 97494 262102
rect 96874 261978 97494 262046
rect 96874 261922 96970 261978
rect 97026 261922 97094 261978
rect 97150 261922 97218 261978
rect 97274 261922 97342 261978
rect 97398 261922 97494 261978
rect 96874 244350 97494 261922
rect 100528 262350 100848 262384
rect 100528 262294 100598 262350
rect 100654 262294 100722 262350
rect 100778 262294 100848 262350
rect 100528 262226 100848 262294
rect 100528 262170 100598 262226
rect 100654 262170 100722 262226
rect 100778 262170 100848 262226
rect 100528 262102 100848 262170
rect 100528 262046 100598 262102
rect 100654 262046 100722 262102
rect 100778 262046 100848 262102
rect 100528 261978 100848 262046
rect 100528 261922 100598 261978
rect 100654 261922 100722 261978
rect 100778 261922 100848 261978
rect 100528 261888 100848 261922
rect 111154 256350 111774 273922
rect 115888 274350 116208 274384
rect 115888 274294 115958 274350
rect 116014 274294 116082 274350
rect 116138 274294 116208 274350
rect 115888 274226 116208 274294
rect 115888 274170 115958 274226
rect 116014 274170 116082 274226
rect 116138 274170 116208 274226
rect 115888 274102 116208 274170
rect 115888 274046 115958 274102
rect 116014 274046 116082 274102
rect 116138 274046 116208 274102
rect 115888 273978 116208 274046
rect 115888 273922 115958 273978
rect 116014 273922 116082 273978
rect 116138 273922 116208 273978
rect 115888 273888 116208 273922
rect 146608 274350 146928 274384
rect 146608 274294 146678 274350
rect 146734 274294 146802 274350
rect 146858 274294 146928 274350
rect 146608 274226 146928 274294
rect 146608 274170 146678 274226
rect 146734 274170 146802 274226
rect 146858 274170 146928 274226
rect 146608 274102 146928 274170
rect 146608 274046 146678 274102
rect 146734 274046 146802 274102
rect 146858 274046 146928 274102
rect 146608 273978 146928 274046
rect 146608 273922 146678 273978
rect 146734 273922 146802 273978
rect 146858 273922 146928 273978
rect 146608 273888 146928 273922
rect 177328 274350 177648 274384
rect 177328 274294 177398 274350
rect 177454 274294 177522 274350
rect 177578 274294 177648 274350
rect 177328 274226 177648 274294
rect 177328 274170 177398 274226
rect 177454 274170 177522 274226
rect 177578 274170 177648 274226
rect 177328 274102 177648 274170
rect 177328 274046 177398 274102
rect 177454 274046 177522 274102
rect 177578 274046 177648 274102
rect 177328 273978 177648 274046
rect 177328 273922 177398 273978
rect 177454 273922 177522 273978
rect 177578 273922 177648 273978
rect 177328 273888 177648 273922
rect 208048 274350 208368 274384
rect 208048 274294 208118 274350
rect 208174 274294 208242 274350
rect 208298 274294 208368 274350
rect 208048 274226 208368 274294
rect 208048 274170 208118 274226
rect 208174 274170 208242 274226
rect 208298 274170 208368 274226
rect 208048 274102 208368 274170
rect 208048 274046 208118 274102
rect 208174 274046 208242 274102
rect 208298 274046 208368 274102
rect 208048 273978 208368 274046
rect 208048 273922 208118 273978
rect 208174 273922 208242 273978
rect 208298 273922 208368 273978
rect 208048 273888 208368 273922
rect 238768 274350 239088 274384
rect 238768 274294 238838 274350
rect 238894 274294 238962 274350
rect 239018 274294 239088 274350
rect 238768 274226 239088 274294
rect 238768 274170 238838 274226
rect 238894 274170 238962 274226
rect 239018 274170 239088 274226
rect 238768 274102 239088 274170
rect 238768 274046 238838 274102
rect 238894 274046 238962 274102
rect 239018 274046 239088 274102
rect 238768 273978 239088 274046
rect 238768 273922 238838 273978
rect 238894 273922 238962 273978
rect 239018 273922 239088 273978
rect 238768 273888 239088 273922
rect 269488 274350 269808 274384
rect 269488 274294 269558 274350
rect 269614 274294 269682 274350
rect 269738 274294 269808 274350
rect 269488 274226 269808 274294
rect 269488 274170 269558 274226
rect 269614 274170 269682 274226
rect 269738 274170 269808 274226
rect 269488 274102 269808 274170
rect 269488 274046 269558 274102
rect 269614 274046 269682 274102
rect 269738 274046 269808 274102
rect 269488 273978 269808 274046
rect 269488 273922 269558 273978
rect 269614 273922 269682 273978
rect 269738 273922 269808 273978
rect 269488 273888 269808 273922
rect 300208 274350 300528 274384
rect 300208 274294 300278 274350
rect 300334 274294 300402 274350
rect 300458 274294 300528 274350
rect 300208 274226 300528 274294
rect 300208 274170 300278 274226
rect 300334 274170 300402 274226
rect 300458 274170 300528 274226
rect 300208 274102 300528 274170
rect 300208 274046 300278 274102
rect 300334 274046 300402 274102
rect 300458 274046 300528 274102
rect 300208 273978 300528 274046
rect 300208 273922 300278 273978
rect 300334 273922 300402 273978
rect 300458 273922 300528 273978
rect 300208 273888 300528 273922
rect 330928 274350 331248 274384
rect 330928 274294 330998 274350
rect 331054 274294 331122 274350
rect 331178 274294 331248 274350
rect 330928 274226 331248 274294
rect 330928 274170 330998 274226
rect 331054 274170 331122 274226
rect 331178 274170 331248 274226
rect 330928 274102 331248 274170
rect 330928 274046 330998 274102
rect 331054 274046 331122 274102
rect 331178 274046 331248 274102
rect 330928 273978 331248 274046
rect 330928 273922 330998 273978
rect 331054 273922 331122 273978
rect 331178 273922 331248 273978
rect 330928 273888 331248 273922
rect 361648 274350 361968 274384
rect 361648 274294 361718 274350
rect 361774 274294 361842 274350
rect 361898 274294 361968 274350
rect 361648 274226 361968 274294
rect 361648 274170 361718 274226
rect 361774 274170 361842 274226
rect 361898 274170 361968 274226
rect 361648 274102 361968 274170
rect 361648 274046 361718 274102
rect 361774 274046 361842 274102
rect 361898 274046 361968 274102
rect 361648 273978 361968 274046
rect 361648 273922 361718 273978
rect 361774 273922 361842 273978
rect 361898 273922 361968 273978
rect 361648 273888 361968 273922
rect 392368 274350 392688 274384
rect 392368 274294 392438 274350
rect 392494 274294 392562 274350
rect 392618 274294 392688 274350
rect 392368 274226 392688 274294
rect 392368 274170 392438 274226
rect 392494 274170 392562 274226
rect 392618 274170 392688 274226
rect 392368 274102 392688 274170
rect 392368 274046 392438 274102
rect 392494 274046 392562 274102
rect 392618 274046 392688 274102
rect 392368 273978 392688 274046
rect 392368 273922 392438 273978
rect 392494 273922 392562 273978
rect 392618 273922 392688 273978
rect 392368 273888 392688 273922
rect 423088 274350 423408 274384
rect 423088 274294 423158 274350
rect 423214 274294 423282 274350
rect 423338 274294 423408 274350
rect 423088 274226 423408 274294
rect 423088 274170 423158 274226
rect 423214 274170 423282 274226
rect 423338 274170 423408 274226
rect 423088 274102 423408 274170
rect 423088 274046 423158 274102
rect 423214 274046 423282 274102
rect 423338 274046 423408 274102
rect 423088 273978 423408 274046
rect 423088 273922 423158 273978
rect 423214 273922 423282 273978
rect 423338 273922 423408 273978
rect 423088 273888 423408 273922
rect 453808 274350 454128 274384
rect 453808 274294 453878 274350
rect 453934 274294 454002 274350
rect 454058 274294 454128 274350
rect 453808 274226 454128 274294
rect 453808 274170 453878 274226
rect 453934 274170 454002 274226
rect 454058 274170 454128 274226
rect 453808 274102 454128 274170
rect 453808 274046 453878 274102
rect 453934 274046 454002 274102
rect 454058 274046 454128 274102
rect 453808 273978 454128 274046
rect 453808 273922 453878 273978
rect 453934 273922 454002 273978
rect 454058 273922 454128 273978
rect 453808 273888 454128 273922
rect 484528 274350 484848 274384
rect 484528 274294 484598 274350
rect 484654 274294 484722 274350
rect 484778 274294 484848 274350
rect 484528 274226 484848 274294
rect 484528 274170 484598 274226
rect 484654 274170 484722 274226
rect 484778 274170 484848 274226
rect 484528 274102 484848 274170
rect 484528 274046 484598 274102
rect 484654 274046 484722 274102
rect 484778 274046 484848 274102
rect 484528 273978 484848 274046
rect 484528 273922 484598 273978
rect 484654 273922 484722 273978
rect 484778 273922 484848 273978
rect 484528 273888 484848 273922
rect 515248 274350 515568 274384
rect 515248 274294 515318 274350
rect 515374 274294 515442 274350
rect 515498 274294 515568 274350
rect 515248 274226 515568 274294
rect 515248 274170 515318 274226
rect 515374 274170 515442 274226
rect 515498 274170 515568 274226
rect 515248 274102 515568 274170
rect 515248 274046 515318 274102
rect 515374 274046 515442 274102
rect 515498 274046 515568 274102
rect 515248 273978 515568 274046
rect 515248 273922 515318 273978
rect 515374 273922 515442 273978
rect 515498 273922 515568 273978
rect 515248 273888 515568 273922
rect 545968 274350 546288 274384
rect 545968 274294 546038 274350
rect 546094 274294 546162 274350
rect 546218 274294 546288 274350
rect 545968 274226 546288 274294
rect 545968 274170 546038 274226
rect 546094 274170 546162 274226
rect 546218 274170 546288 274226
rect 545968 274102 546288 274170
rect 545968 274046 546038 274102
rect 546094 274046 546162 274102
rect 546218 274046 546288 274102
rect 545968 273978 546288 274046
rect 545968 273922 546038 273978
rect 546094 273922 546162 273978
rect 546218 273922 546288 273978
rect 545968 273888 546288 273922
rect 561154 274350 561774 291922
rect 561154 274294 561250 274350
rect 561306 274294 561374 274350
rect 561430 274294 561498 274350
rect 561554 274294 561622 274350
rect 561678 274294 561774 274350
rect 561154 274226 561774 274294
rect 561154 274170 561250 274226
rect 561306 274170 561374 274226
rect 561430 274170 561498 274226
rect 561554 274170 561622 274226
rect 561678 274170 561774 274226
rect 561154 274102 561774 274170
rect 561154 274046 561250 274102
rect 561306 274046 561374 274102
rect 561430 274046 561498 274102
rect 561554 274046 561622 274102
rect 561678 274046 561774 274102
rect 561154 273978 561774 274046
rect 561154 273922 561250 273978
rect 561306 273922 561374 273978
rect 561430 273922 561498 273978
rect 561554 273922 561622 273978
rect 561678 273922 561774 273978
rect 131248 262350 131568 262384
rect 131248 262294 131318 262350
rect 131374 262294 131442 262350
rect 131498 262294 131568 262350
rect 131248 262226 131568 262294
rect 131248 262170 131318 262226
rect 131374 262170 131442 262226
rect 131498 262170 131568 262226
rect 131248 262102 131568 262170
rect 131248 262046 131318 262102
rect 131374 262046 131442 262102
rect 131498 262046 131568 262102
rect 131248 261978 131568 262046
rect 131248 261922 131318 261978
rect 131374 261922 131442 261978
rect 131498 261922 131568 261978
rect 131248 261888 131568 261922
rect 161968 262350 162288 262384
rect 161968 262294 162038 262350
rect 162094 262294 162162 262350
rect 162218 262294 162288 262350
rect 161968 262226 162288 262294
rect 161968 262170 162038 262226
rect 162094 262170 162162 262226
rect 162218 262170 162288 262226
rect 161968 262102 162288 262170
rect 161968 262046 162038 262102
rect 162094 262046 162162 262102
rect 162218 262046 162288 262102
rect 161968 261978 162288 262046
rect 161968 261922 162038 261978
rect 162094 261922 162162 261978
rect 162218 261922 162288 261978
rect 161968 261888 162288 261922
rect 192688 262350 193008 262384
rect 192688 262294 192758 262350
rect 192814 262294 192882 262350
rect 192938 262294 193008 262350
rect 192688 262226 193008 262294
rect 192688 262170 192758 262226
rect 192814 262170 192882 262226
rect 192938 262170 193008 262226
rect 192688 262102 193008 262170
rect 192688 262046 192758 262102
rect 192814 262046 192882 262102
rect 192938 262046 193008 262102
rect 192688 261978 193008 262046
rect 192688 261922 192758 261978
rect 192814 261922 192882 261978
rect 192938 261922 193008 261978
rect 192688 261888 193008 261922
rect 223408 262350 223728 262384
rect 223408 262294 223478 262350
rect 223534 262294 223602 262350
rect 223658 262294 223728 262350
rect 223408 262226 223728 262294
rect 223408 262170 223478 262226
rect 223534 262170 223602 262226
rect 223658 262170 223728 262226
rect 223408 262102 223728 262170
rect 223408 262046 223478 262102
rect 223534 262046 223602 262102
rect 223658 262046 223728 262102
rect 223408 261978 223728 262046
rect 223408 261922 223478 261978
rect 223534 261922 223602 261978
rect 223658 261922 223728 261978
rect 223408 261888 223728 261922
rect 254128 262350 254448 262384
rect 254128 262294 254198 262350
rect 254254 262294 254322 262350
rect 254378 262294 254448 262350
rect 254128 262226 254448 262294
rect 254128 262170 254198 262226
rect 254254 262170 254322 262226
rect 254378 262170 254448 262226
rect 254128 262102 254448 262170
rect 254128 262046 254198 262102
rect 254254 262046 254322 262102
rect 254378 262046 254448 262102
rect 254128 261978 254448 262046
rect 254128 261922 254198 261978
rect 254254 261922 254322 261978
rect 254378 261922 254448 261978
rect 254128 261888 254448 261922
rect 284848 262350 285168 262384
rect 284848 262294 284918 262350
rect 284974 262294 285042 262350
rect 285098 262294 285168 262350
rect 284848 262226 285168 262294
rect 284848 262170 284918 262226
rect 284974 262170 285042 262226
rect 285098 262170 285168 262226
rect 284848 262102 285168 262170
rect 284848 262046 284918 262102
rect 284974 262046 285042 262102
rect 285098 262046 285168 262102
rect 284848 261978 285168 262046
rect 284848 261922 284918 261978
rect 284974 261922 285042 261978
rect 285098 261922 285168 261978
rect 284848 261888 285168 261922
rect 315568 262350 315888 262384
rect 315568 262294 315638 262350
rect 315694 262294 315762 262350
rect 315818 262294 315888 262350
rect 315568 262226 315888 262294
rect 315568 262170 315638 262226
rect 315694 262170 315762 262226
rect 315818 262170 315888 262226
rect 315568 262102 315888 262170
rect 315568 262046 315638 262102
rect 315694 262046 315762 262102
rect 315818 262046 315888 262102
rect 315568 261978 315888 262046
rect 315568 261922 315638 261978
rect 315694 261922 315762 261978
rect 315818 261922 315888 261978
rect 315568 261888 315888 261922
rect 346288 262350 346608 262384
rect 346288 262294 346358 262350
rect 346414 262294 346482 262350
rect 346538 262294 346608 262350
rect 346288 262226 346608 262294
rect 346288 262170 346358 262226
rect 346414 262170 346482 262226
rect 346538 262170 346608 262226
rect 346288 262102 346608 262170
rect 346288 262046 346358 262102
rect 346414 262046 346482 262102
rect 346538 262046 346608 262102
rect 346288 261978 346608 262046
rect 346288 261922 346358 261978
rect 346414 261922 346482 261978
rect 346538 261922 346608 261978
rect 346288 261888 346608 261922
rect 377008 262350 377328 262384
rect 377008 262294 377078 262350
rect 377134 262294 377202 262350
rect 377258 262294 377328 262350
rect 377008 262226 377328 262294
rect 377008 262170 377078 262226
rect 377134 262170 377202 262226
rect 377258 262170 377328 262226
rect 377008 262102 377328 262170
rect 377008 262046 377078 262102
rect 377134 262046 377202 262102
rect 377258 262046 377328 262102
rect 377008 261978 377328 262046
rect 377008 261922 377078 261978
rect 377134 261922 377202 261978
rect 377258 261922 377328 261978
rect 377008 261888 377328 261922
rect 407728 262350 408048 262384
rect 407728 262294 407798 262350
rect 407854 262294 407922 262350
rect 407978 262294 408048 262350
rect 407728 262226 408048 262294
rect 407728 262170 407798 262226
rect 407854 262170 407922 262226
rect 407978 262170 408048 262226
rect 407728 262102 408048 262170
rect 407728 262046 407798 262102
rect 407854 262046 407922 262102
rect 407978 262046 408048 262102
rect 407728 261978 408048 262046
rect 407728 261922 407798 261978
rect 407854 261922 407922 261978
rect 407978 261922 408048 261978
rect 407728 261888 408048 261922
rect 438448 262350 438768 262384
rect 438448 262294 438518 262350
rect 438574 262294 438642 262350
rect 438698 262294 438768 262350
rect 438448 262226 438768 262294
rect 438448 262170 438518 262226
rect 438574 262170 438642 262226
rect 438698 262170 438768 262226
rect 438448 262102 438768 262170
rect 438448 262046 438518 262102
rect 438574 262046 438642 262102
rect 438698 262046 438768 262102
rect 438448 261978 438768 262046
rect 438448 261922 438518 261978
rect 438574 261922 438642 261978
rect 438698 261922 438768 261978
rect 438448 261888 438768 261922
rect 469168 262350 469488 262384
rect 469168 262294 469238 262350
rect 469294 262294 469362 262350
rect 469418 262294 469488 262350
rect 469168 262226 469488 262294
rect 469168 262170 469238 262226
rect 469294 262170 469362 262226
rect 469418 262170 469488 262226
rect 469168 262102 469488 262170
rect 469168 262046 469238 262102
rect 469294 262046 469362 262102
rect 469418 262046 469488 262102
rect 469168 261978 469488 262046
rect 469168 261922 469238 261978
rect 469294 261922 469362 261978
rect 469418 261922 469488 261978
rect 469168 261888 469488 261922
rect 499888 262350 500208 262384
rect 499888 262294 499958 262350
rect 500014 262294 500082 262350
rect 500138 262294 500208 262350
rect 499888 262226 500208 262294
rect 499888 262170 499958 262226
rect 500014 262170 500082 262226
rect 500138 262170 500208 262226
rect 499888 262102 500208 262170
rect 499888 262046 499958 262102
rect 500014 262046 500082 262102
rect 500138 262046 500208 262102
rect 499888 261978 500208 262046
rect 499888 261922 499958 261978
rect 500014 261922 500082 261978
rect 500138 261922 500208 261978
rect 499888 261888 500208 261922
rect 530608 262350 530928 262384
rect 530608 262294 530678 262350
rect 530734 262294 530802 262350
rect 530858 262294 530928 262350
rect 530608 262226 530928 262294
rect 530608 262170 530678 262226
rect 530734 262170 530802 262226
rect 530858 262170 530928 262226
rect 530608 262102 530928 262170
rect 530608 262046 530678 262102
rect 530734 262046 530802 262102
rect 530858 262046 530928 262102
rect 530608 261978 530928 262046
rect 530608 261922 530678 261978
rect 530734 261922 530802 261978
rect 530858 261922 530928 261978
rect 530608 261888 530928 261922
rect 111154 256294 111250 256350
rect 111306 256294 111374 256350
rect 111430 256294 111498 256350
rect 111554 256294 111622 256350
rect 111678 256294 111774 256350
rect 111154 256226 111774 256294
rect 111154 256170 111250 256226
rect 111306 256170 111374 256226
rect 111430 256170 111498 256226
rect 111554 256170 111622 256226
rect 111678 256170 111774 256226
rect 111154 256102 111774 256170
rect 111154 256046 111250 256102
rect 111306 256046 111374 256102
rect 111430 256046 111498 256102
rect 111554 256046 111622 256102
rect 111678 256046 111774 256102
rect 111154 255978 111774 256046
rect 111154 255922 111250 255978
rect 111306 255922 111374 255978
rect 111430 255922 111498 255978
rect 111554 255922 111622 255978
rect 111678 255922 111774 255978
rect 96874 244294 96970 244350
rect 97026 244294 97094 244350
rect 97150 244294 97218 244350
rect 97274 244294 97342 244350
rect 97398 244294 97494 244350
rect 96874 244226 97494 244294
rect 96874 244170 96970 244226
rect 97026 244170 97094 244226
rect 97150 244170 97218 244226
rect 97274 244170 97342 244226
rect 97398 244170 97494 244226
rect 96874 244102 97494 244170
rect 96874 244046 96970 244102
rect 97026 244046 97094 244102
rect 97150 244046 97218 244102
rect 97274 244046 97342 244102
rect 97398 244046 97494 244102
rect 96874 243978 97494 244046
rect 96874 243922 96970 243978
rect 97026 243922 97094 243978
rect 97150 243922 97218 243978
rect 97274 243922 97342 243978
rect 97398 243922 97494 243978
rect 96874 226350 97494 243922
rect 100528 244350 100848 244384
rect 100528 244294 100598 244350
rect 100654 244294 100722 244350
rect 100778 244294 100848 244350
rect 100528 244226 100848 244294
rect 100528 244170 100598 244226
rect 100654 244170 100722 244226
rect 100778 244170 100848 244226
rect 100528 244102 100848 244170
rect 100528 244046 100598 244102
rect 100654 244046 100722 244102
rect 100778 244046 100848 244102
rect 100528 243978 100848 244046
rect 100528 243922 100598 243978
rect 100654 243922 100722 243978
rect 100778 243922 100848 243978
rect 100528 243888 100848 243922
rect 111154 238350 111774 255922
rect 115888 256350 116208 256384
rect 115888 256294 115958 256350
rect 116014 256294 116082 256350
rect 116138 256294 116208 256350
rect 115888 256226 116208 256294
rect 115888 256170 115958 256226
rect 116014 256170 116082 256226
rect 116138 256170 116208 256226
rect 115888 256102 116208 256170
rect 115888 256046 115958 256102
rect 116014 256046 116082 256102
rect 116138 256046 116208 256102
rect 115888 255978 116208 256046
rect 115888 255922 115958 255978
rect 116014 255922 116082 255978
rect 116138 255922 116208 255978
rect 115888 255888 116208 255922
rect 146608 256350 146928 256384
rect 146608 256294 146678 256350
rect 146734 256294 146802 256350
rect 146858 256294 146928 256350
rect 146608 256226 146928 256294
rect 146608 256170 146678 256226
rect 146734 256170 146802 256226
rect 146858 256170 146928 256226
rect 146608 256102 146928 256170
rect 146608 256046 146678 256102
rect 146734 256046 146802 256102
rect 146858 256046 146928 256102
rect 146608 255978 146928 256046
rect 146608 255922 146678 255978
rect 146734 255922 146802 255978
rect 146858 255922 146928 255978
rect 146608 255888 146928 255922
rect 177328 256350 177648 256384
rect 177328 256294 177398 256350
rect 177454 256294 177522 256350
rect 177578 256294 177648 256350
rect 177328 256226 177648 256294
rect 177328 256170 177398 256226
rect 177454 256170 177522 256226
rect 177578 256170 177648 256226
rect 177328 256102 177648 256170
rect 177328 256046 177398 256102
rect 177454 256046 177522 256102
rect 177578 256046 177648 256102
rect 177328 255978 177648 256046
rect 177328 255922 177398 255978
rect 177454 255922 177522 255978
rect 177578 255922 177648 255978
rect 177328 255888 177648 255922
rect 208048 256350 208368 256384
rect 208048 256294 208118 256350
rect 208174 256294 208242 256350
rect 208298 256294 208368 256350
rect 208048 256226 208368 256294
rect 208048 256170 208118 256226
rect 208174 256170 208242 256226
rect 208298 256170 208368 256226
rect 208048 256102 208368 256170
rect 208048 256046 208118 256102
rect 208174 256046 208242 256102
rect 208298 256046 208368 256102
rect 208048 255978 208368 256046
rect 208048 255922 208118 255978
rect 208174 255922 208242 255978
rect 208298 255922 208368 255978
rect 208048 255888 208368 255922
rect 238768 256350 239088 256384
rect 238768 256294 238838 256350
rect 238894 256294 238962 256350
rect 239018 256294 239088 256350
rect 238768 256226 239088 256294
rect 238768 256170 238838 256226
rect 238894 256170 238962 256226
rect 239018 256170 239088 256226
rect 238768 256102 239088 256170
rect 238768 256046 238838 256102
rect 238894 256046 238962 256102
rect 239018 256046 239088 256102
rect 238768 255978 239088 256046
rect 238768 255922 238838 255978
rect 238894 255922 238962 255978
rect 239018 255922 239088 255978
rect 238768 255888 239088 255922
rect 269488 256350 269808 256384
rect 269488 256294 269558 256350
rect 269614 256294 269682 256350
rect 269738 256294 269808 256350
rect 269488 256226 269808 256294
rect 269488 256170 269558 256226
rect 269614 256170 269682 256226
rect 269738 256170 269808 256226
rect 269488 256102 269808 256170
rect 269488 256046 269558 256102
rect 269614 256046 269682 256102
rect 269738 256046 269808 256102
rect 269488 255978 269808 256046
rect 269488 255922 269558 255978
rect 269614 255922 269682 255978
rect 269738 255922 269808 255978
rect 269488 255888 269808 255922
rect 300208 256350 300528 256384
rect 300208 256294 300278 256350
rect 300334 256294 300402 256350
rect 300458 256294 300528 256350
rect 300208 256226 300528 256294
rect 300208 256170 300278 256226
rect 300334 256170 300402 256226
rect 300458 256170 300528 256226
rect 300208 256102 300528 256170
rect 300208 256046 300278 256102
rect 300334 256046 300402 256102
rect 300458 256046 300528 256102
rect 300208 255978 300528 256046
rect 300208 255922 300278 255978
rect 300334 255922 300402 255978
rect 300458 255922 300528 255978
rect 300208 255888 300528 255922
rect 330928 256350 331248 256384
rect 330928 256294 330998 256350
rect 331054 256294 331122 256350
rect 331178 256294 331248 256350
rect 330928 256226 331248 256294
rect 330928 256170 330998 256226
rect 331054 256170 331122 256226
rect 331178 256170 331248 256226
rect 330928 256102 331248 256170
rect 330928 256046 330998 256102
rect 331054 256046 331122 256102
rect 331178 256046 331248 256102
rect 330928 255978 331248 256046
rect 330928 255922 330998 255978
rect 331054 255922 331122 255978
rect 331178 255922 331248 255978
rect 330928 255888 331248 255922
rect 361648 256350 361968 256384
rect 361648 256294 361718 256350
rect 361774 256294 361842 256350
rect 361898 256294 361968 256350
rect 361648 256226 361968 256294
rect 361648 256170 361718 256226
rect 361774 256170 361842 256226
rect 361898 256170 361968 256226
rect 361648 256102 361968 256170
rect 361648 256046 361718 256102
rect 361774 256046 361842 256102
rect 361898 256046 361968 256102
rect 361648 255978 361968 256046
rect 361648 255922 361718 255978
rect 361774 255922 361842 255978
rect 361898 255922 361968 255978
rect 361648 255888 361968 255922
rect 392368 256350 392688 256384
rect 392368 256294 392438 256350
rect 392494 256294 392562 256350
rect 392618 256294 392688 256350
rect 392368 256226 392688 256294
rect 392368 256170 392438 256226
rect 392494 256170 392562 256226
rect 392618 256170 392688 256226
rect 392368 256102 392688 256170
rect 392368 256046 392438 256102
rect 392494 256046 392562 256102
rect 392618 256046 392688 256102
rect 392368 255978 392688 256046
rect 392368 255922 392438 255978
rect 392494 255922 392562 255978
rect 392618 255922 392688 255978
rect 392368 255888 392688 255922
rect 423088 256350 423408 256384
rect 423088 256294 423158 256350
rect 423214 256294 423282 256350
rect 423338 256294 423408 256350
rect 423088 256226 423408 256294
rect 423088 256170 423158 256226
rect 423214 256170 423282 256226
rect 423338 256170 423408 256226
rect 423088 256102 423408 256170
rect 423088 256046 423158 256102
rect 423214 256046 423282 256102
rect 423338 256046 423408 256102
rect 423088 255978 423408 256046
rect 423088 255922 423158 255978
rect 423214 255922 423282 255978
rect 423338 255922 423408 255978
rect 423088 255888 423408 255922
rect 453808 256350 454128 256384
rect 453808 256294 453878 256350
rect 453934 256294 454002 256350
rect 454058 256294 454128 256350
rect 453808 256226 454128 256294
rect 453808 256170 453878 256226
rect 453934 256170 454002 256226
rect 454058 256170 454128 256226
rect 453808 256102 454128 256170
rect 453808 256046 453878 256102
rect 453934 256046 454002 256102
rect 454058 256046 454128 256102
rect 453808 255978 454128 256046
rect 453808 255922 453878 255978
rect 453934 255922 454002 255978
rect 454058 255922 454128 255978
rect 453808 255888 454128 255922
rect 484528 256350 484848 256384
rect 484528 256294 484598 256350
rect 484654 256294 484722 256350
rect 484778 256294 484848 256350
rect 484528 256226 484848 256294
rect 484528 256170 484598 256226
rect 484654 256170 484722 256226
rect 484778 256170 484848 256226
rect 484528 256102 484848 256170
rect 484528 256046 484598 256102
rect 484654 256046 484722 256102
rect 484778 256046 484848 256102
rect 484528 255978 484848 256046
rect 484528 255922 484598 255978
rect 484654 255922 484722 255978
rect 484778 255922 484848 255978
rect 484528 255888 484848 255922
rect 515248 256350 515568 256384
rect 515248 256294 515318 256350
rect 515374 256294 515442 256350
rect 515498 256294 515568 256350
rect 515248 256226 515568 256294
rect 515248 256170 515318 256226
rect 515374 256170 515442 256226
rect 515498 256170 515568 256226
rect 515248 256102 515568 256170
rect 515248 256046 515318 256102
rect 515374 256046 515442 256102
rect 515498 256046 515568 256102
rect 515248 255978 515568 256046
rect 515248 255922 515318 255978
rect 515374 255922 515442 255978
rect 515498 255922 515568 255978
rect 515248 255888 515568 255922
rect 545968 256350 546288 256384
rect 545968 256294 546038 256350
rect 546094 256294 546162 256350
rect 546218 256294 546288 256350
rect 545968 256226 546288 256294
rect 545968 256170 546038 256226
rect 546094 256170 546162 256226
rect 546218 256170 546288 256226
rect 545968 256102 546288 256170
rect 545968 256046 546038 256102
rect 546094 256046 546162 256102
rect 546218 256046 546288 256102
rect 545968 255978 546288 256046
rect 545968 255922 546038 255978
rect 546094 255922 546162 255978
rect 546218 255922 546288 255978
rect 545968 255888 546288 255922
rect 561154 256350 561774 273922
rect 561154 256294 561250 256350
rect 561306 256294 561374 256350
rect 561430 256294 561498 256350
rect 561554 256294 561622 256350
rect 561678 256294 561774 256350
rect 561154 256226 561774 256294
rect 561154 256170 561250 256226
rect 561306 256170 561374 256226
rect 561430 256170 561498 256226
rect 561554 256170 561622 256226
rect 561678 256170 561774 256226
rect 561154 256102 561774 256170
rect 561154 256046 561250 256102
rect 561306 256046 561374 256102
rect 561430 256046 561498 256102
rect 561554 256046 561622 256102
rect 561678 256046 561774 256102
rect 561154 255978 561774 256046
rect 561154 255922 561250 255978
rect 561306 255922 561374 255978
rect 561430 255922 561498 255978
rect 561554 255922 561622 255978
rect 561678 255922 561774 255978
rect 131248 244350 131568 244384
rect 131248 244294 131318 244350
rect 131374 244294 131442 244350
rect 131498 244294 131568 244350
rect 131248 244226 131568 244294
rect 131248 244170 131318 244226
rect 131374 244170 131442 244226
rect 131498 244170 131568 244226
rect 131248 244102 131568 244170
rect 131248 244046 131318 244102
rect 131374 244046 131442 244102
rect 131498 244046 131568 244102
rect 131248 243978 131568 244046
rect 131248 243922 131318 243978
rect 131374 243922 131442 243978
rect 131498 243922 131568 243978
rect 131248 243888 131568 243922
rect 161968 244350 162288 244384
rect 161968 244294 162038 244350
rect 162094 244294 162162 244350
rect 162218 244294 162288 244350
rect 161968 244226 162288 244294
rect 161968 244170 162038 244226
rect 162094 244170 162162 244226
rect 162218 244170 162288 244226
rect 161968 244102 162288 244170
rect 161968 244046 162038 244102
rect 162094 244046 162162 244102
rect 162218 244046 162288 244102
rect 161968 243978 162288 244046
rect 161968 243922 162038 243978
rect 162094 243922 162162 243978
rect 162218 243922 162288 243978
rect 161968 243888 162288 243922
rect 192688 244350 193008 244384
rect 192688 244294 192758 244350
rect 192814 244294 192882 244350
rect 192938 244294 193008 244350
rect 192688 244226 193008 244294
rect 192688 244170 192758 244226
rect 192814 244170 192882 244226
rect 192938 244170 193008 244226
rect 192688 244102 193008 244170
rect 192688 244046 192758 244102
rect 192814 244046 192882 244102
rect 192938 244046 193008 244102
rect 192688 243978 193008 244046
rect 192688 243922 192758 243978
rect 192814 243922 192882 243978
rect 192938 243922 193008 243978
rect 192688 243888 193008 243922
rect 223408 244350 223728 244384
rect 223408 244294 223478 244350
rect 223534 244294 223602 244350
rect 223658 244294 223728 244350
rect 223408 244226 223728 244294
rect 223408 244170 223478 244226
rect 223534 244170 223602 244226
rect 223658 244170 223728 244226
rect 223408 244102 223728 244170
rect 223408 244046 223478 244102
rect 223534 244046 223602 244102
rect 223658 244046 223728 244102
rect 223408 243978 223728 244046
rect 223408 243922 223478 243978
rect 223534 243922 223602 243978
rect 223658 243922 223728 243978
rect 223408 243888 223728 243922
rect 254128 244350 254448 244384
rect 254128 244294 254198 244350
rect 254254 244294 254322 244350
rect 254378 244294 254448 244350
rect 254128 244226 254448 244294
rect 254128 244170 254198 244226
rect 254254 244170 254322 244226
rect 254378 244170 254448 244226
rect 254128 244102 254448 244170
rect 254128 244046 254198 244102
rect 254254 244046 254322 244102
rect 254378 244046 254448 244102
rect 254128 243978 254448 244046
rect 254128 243922 254198 243978
rect 254254 243922 254322 243978
rect 254378 243922 254448 243978
rect 254128 243888 254448 243922
rect 284848 244350 285168 244384
rect 284848 244294 284918 244350
rect 284974 244294 285042 244350
rect 285098 244294 285168 244350
rect 284848 244226 285168 244294
rect 284848 244170 284918 244226
rect 284974 244170 285042 244226
rect 285098 244170 285168 244226
rect 284848 244102 285168 244170
rect 284848 244046 284918 244102
rect 284974 244046 285042 244102
rect 285098 244046 285168 244102
rect 284848 243978 285168 244046
rect 284848 243922 284918 243978
rect 284974 243922 285042 243978
rect 285098 243922 285168 243978
rect 284848 243888 285168 243922
rect 315568 244350 315888 244384
rect 315568 244294 315638 244350
rect 315694 244294 315762 244350
rect 315818 244294 315888 244350
rect 315568 244226 315888 244294
rect 315568 244170 315638 244226
rect 315694 244170 315762 244226
rect 315818 244170 315888 244226
rect 315568 244102 315888 244170
rect 315568 244046 315638 244102
rect 315694 244046 315762 244102
rect 315818 244046 315888 244102
rect 315568 243978 315888 244046
rect 315568 243922 315638 243978
rect 315694 243922 315762 243978
rect 315818 243922 315888 243978
rect 315568 243888 315888 243922
rect 346288 244350 346608 244384
rect 346288 244294 346358 244350
rect 346414 244294 346482 244350
rect 346538 244294 346608 244350
rect 346288 244226 346608 244294
rect 346288 244170 346358 244226
rect 346414 244170 346482 244226
rect 346538 244170 346608 244226
rect 346288 244102 346608 244170
rect 346288 244046 346358 244102
rect 346414 244046 346482 244102
rect 346538 244046 346608 244102
rect 346288 243978 346608 244046
rect 346288 243922 346358 243978
rect 346414 243922 346482 243978
rect 346538 243922 346608 243978
rect 346288 243888 346608 243922
rect 377008 244350 377328 244384
rect 377008 244294 377078 244350
rect 377134 244294 377202 244350
rect 377258 244294 377328 244350
rect 377008 244226 377328 244294
rect 377008 244170 377078 244226
rect 377134 244170 377202 244226
rect 377258 244170 377328 244226
rect 377008 244102 377328 244170
rect 377008 244046 377078 244102
rect 377134 244046 377202 244102
rect 377258 244046 377328 244102
rect 377008 243978 377328 244046
rect 377008 243922 377078 243978
rect 377134 243922 377202 243978
rect 377258 243922 377328 243978
rect 377008 243888 377328 243922
rect 407728 244350 408048 244384
rect 407728 244294 407798 244350
rect 407854 244294 407922 244350
rect 407978 244294 408048 244350
rect 407728 244226 408048 244294
rect 407728 244170 407798 244226
rect 407854 244170 407922 244226
rect 407978 244170 408048 244226
rect 407728 244102 408048 244170
rect 407728 244046 407798 244102
rect 407854 244046 407922 244102
rect 407978 244046 408048 244102
rect 407728 243978 408048 244046
rect 407728 243922 407798 243978
rect 407854 243922 407922 243978
rect 407978 243922 408048 243978
rect 407728 243888 408048 243922
rect 438448 244350 438768 244384
rect 438448 244294 438518 244350
rect 438574 244294 438642 244350
rect 438698 244294 438768 244350
rect 438448 244226 438768 244294
rect 438448 244170 438518 244226
rect 438574 244170 438642 244226
rect 438698 244170 438768 244226
rect 438448 244102 438768 244170
rect 438448 244046 438518 244102
rect 438574 244046 438642 244102
rect 438698 244046 438768 244102
rect 438448 243978 438768 244046
rect 438448 243922 438518 243978
rect 438574 243922 438642 243978
rect 438698 243922 438768 243978
rect 438448 243888 438768 243922
rect 469168 244350 469488 244384
rect 469168 244294 469238 244350
rect 469294 244294 469362 244350
rect 469418 244294 469488 244350
rect 469168 244226 469488 244294
rect 469168 244170 469238 244226
rect 469294 244170 469362 244226
rect 469418 244170 469488 244226
rect 469168 244102 469488 244170
rect 469168 244046 469238 244102
rect 469294 244046 469362 244102
rect 469418 244046 469488 244102
rect 469168 243978 469488 244046
rect 469168 243922 469238 243978
rect 469294 243922 469362 243978
rect 469418 243922 469488 243978
rect 469168 243888 469488 243922
rect 499888 244350 500208 244384
rect 499888 244294 499958 244350
rect 500014 244294 500082 244350
rect 500138 244294 500208 244350
rect 499888 244226 500208 244294
rect 499888 244170 499958 244226
rect 500014 244170 500082 244226
rect 500138 244170 500208 244226
rect 499888 244102 500208 244170
rect 499888 244046 499958 244102
rect 500014 244046 500082 244102
rect 500138 244046 500208 244102
rect 499888 243978 500208 244046
rect 499888 243922 499958 243978
rect 500014 243922 500082 243978
rect 500138 243922 500208 243978
rect 499888 243888 500208 243922
rect 530608 244350 530928 244384
rect 530608 244294 530678 244350
rect 530734 244294 530802 244350
rect 530858 244294 530928 244350
rect 530608 244226 530928 244294
rect 530608 244170 530678 244226
rect 530734 244170 530802 244226
rect 530858 244170 530928 244226
rect 530608 244102 530928 244170
rect 530608 244046 530678 244102
rect 530734 244046 530802 244102
rect 530858 244046 530928 244102
rect 530608 243978 530928 244046
rect 530608 243922 530678 243978
rect 530734 243922 530802 243978
rect 530858 243922 530928 243978
rect 530608 243888 530928 243922
rect 111154 238294 111250 238350
rect 111306 238294 111374 238350
rect 111430 238294 111498 238350
rect 111554 238294 111622 238350
rect 111678 238294 111774 238350
rect 111154 238226 111774 238294
rect 111154 238170 111250 238226
rect 111306 238170 111374 238226
rect 111430 238170 111498 238226
rect 111554 238170 111622 238226
rect 111678 238170 111774 238226
rect 111154 238102 111774 238170
rect 111154 238046 111250 238102
rect 111306 238046 111374 238102
rect 111430 238046 111498 238102
rect 111554 238046 111622 238102
rect 111678 238046 111774 238102
rect 111154 237978 111774 238046
rect 111154 237922 111250 237978
rect 111306 237922 111374 237978
rect 111430 237922 111498 237978
rect 111554 237922 111622 237978
rect 111678 237922 111774 237978
rect 96874 226294 96970 226350
rect 97026 226294 97094 226350
rect 97150 226294 97218 226350
rect 97274 226294 97342 226350
rect 97398 226294 97494 226350
rect 96874 226226 97494 226294
rect 96874 226170 96970 226226
rect 97026 226170 97094 226226
rect 97150 226170 97218 226226
rect 97274 226170 97342 226226
rect 97398 226170 97494 226226
rect 96874 226102 97494 226170
rect 96874 226046 96970 226102
rect 97026 226046 97094 226102
rect 97150 226046 97218 226102
rect 97274 226046 97342 226102
rect 97398 226046 97494 226102
rect 96874 225978 97494 226046
rect 96874 225922 96970 225978
rect 97026 225922 97094 225978
rect 97150 225922 97218 225978
rect 97274 225922 97342 225978
rect 97398 225922 97494 225978
rect 96874 208350 97494 225922
rect 100528 226350 100848 226384
rect 100528 226294 100598 226350
rect 100654 226294 100722 226350
rect 100778 226294 100848 226350
rect 100528 226226 100848 226294
rect 100528 226170 100598 226226
rect 100654 226170 100722 226226
rect 100778 226170 100848 226226
rect 100528 226102 100848 226170
rect 100528 226046 100598 226102
rect 100654 226046 100722 226102
rect 100778 226046 100848 226102
rect 100528 225978 100848 226046
rect 100528 225922 100598 225978
rect 100654 225922 100722 225978
rect 100778 225922 100848 225978
rect 100528 225888 100848 225922
rect 111154 220350 111774 237922
rect 115888 238350 116208 238384
rect 115888 238294 115958 238350
rect 116014 238294 116082 238350
rect 116138 238294 116208 238350
rect 115888 238226 116208 238294
rect 115888 238170 115958 238226
rect 116014 238170 116082 238226
rect 116138 238170 116208 238226
rect 115888 238102 116208 238170
rect 115888 238046 115958 238102
rect 116014 238046 116082 238102
rect 116138 238046 116208 238102
rect 115888 237978 116208 238046
rect 115888 237922 115958 237978
rect 116014 237922 116082 237978
rect 116138 237922 116208 237978
rect 115888 237888 116208 237922
rect 146608 238350 146928 238384
rect 146608 238294 146678 238350
rect 146734 238294 146802 238350
rect 146858 238294 146928 238350
rect 146608 238226 146928 238294
rect 146608 238170 146678 238226
rect 146734 238170 146802 238226
rect 146858 238170 146928 238226
rect 146608 238102 146928 238170
rect 146608 238046 146678 238102
rect 146734 238046 146802 238102
rect 146858 238046 146928 238102
rect 146608 237978 146928 238046
rect 146608 237922 146678 237978
rect 146734 237922 146802 237978
rect 146858 237922 146928 237978
rect 146608 237888 146928 237922
rect 177328 238350 177648 238384
rect 177328 238294 177398 238350
rect 177454 238294 177522 238350
rect 177578 238294 177648 238350
rect 177328 238226 177648 238294
rect 177328 238170 177398 238226
rect 177454 238170 177522 238226
rect 177578 238170 177648 238226
rect 177328 238102 177648 238170
rect 177328 238046 177398 238102
rect 177454 238046 177522 238102
rect 177578 238046 177648 238102
rect 177328 237978 177648 238046
rect 177328 237922 177398 237978
rect 177454 237922 177522 237978
rect 177578 237922 177648 237978
rect 177328 237888 177648 237922
rect 208048 238350 208368 238384
rect 208048 238294 208118 238350
rect 208174 238294 208242 238350
rect 208298 238294 208368 238350
rect 208048 238226 208368 238294
rect 208048 238170 208118 238226
rect 208174 238170 208242 238226
rect 208298 238170 208368 238226
rect 208048 238102 208368 238170
rect 208048 238046 208118 238102
rect 208174 238046 208242 238102
rect 208298 238046 208368 238102
rect 208048 237978 208368 238046
rect 208048 237922 208118 237978
rect 208174 237922 208242 237978
rect 208298 237922 208368 237978
rect 208048 237888 208368 237922
rect 238768 238350 239088 238384
rect 238768 238294 238838 238350
rect 238894 238294 238962 238350
rect 239018 238294 239088 238350
rect 238768 238226 239088 238294
rect 238768 238170 238838 238226
rect 238894 238170 238962 238226
rect 239018 238170 239088 238226
rect 238768 238102 239088 238170
rect 238768 238046 238838 238102
rect 238894 238046 238962 238102
rect 239018 238046 239088 238102
rect 238768 237978 239088 238046
rect 238768 237922 238838 237978
rect 238894 237922 238962 237978
rect 239018 237922 239088 237978
rect 238768 237888 239088 237922
rect 269488 238350 269808 238384
rect 269488 238294 269558 238350
rect 269614 238294 269682 238350
rect 269738 238294 269808 238350
rect 269488 238226 269808 238294
rect 269488 238170 269558 238226
rect 269614 238170 269682 238226
rect 269738 238170 269808 238226
rect 269488 238102 269808 238170
rect 269488 238046 269558 238102
rect 269614 238046 269682 238102
rect 269738 238046 269808 238102
rect 269488 237978 269808 238046
rect 269488 237922 269558 237978
rect 269614 237922 269682 237978
rect 269738 237922 269808 237978
rect 269488 237888 269808 237922
rect 300208 238350 300528 238384
rect 300208 238294 300278 238350
rect 300334 238294 300402 238350
rect 300458 238294 300528 238350
rect 300208 238226 300528 238294
rect 300208 238170 300278 238226
rect 300334 238170 300402 238226
rect 300458 238170 300528 238226
rect 300208 238102 300528 238170
rect 300208 238046 300278 238102
rect 300334 238046 300402 238102
rect 300458 238046 300528 238102
rect 300208 237978 300528 238046
rect 300208 237922 300278 237978
rect 300334 237922 300402 237978
rect 300458 237922 300528 237978
rect 300208 237888 300528 237922
rect 330928 238350 331248 238384
rect 330928 238294 330998 238350
rect 331054 238294 331122 238350
rect 331178 238294 331248 238350
rect 330928 238226 331248 238294
rect 330928 238170 330998 238226
rect 331054 238170 331122 238226
rect 331178 238170 331248 238226
rect 330928 238102 331248 238170
rect 330928 238046 330998 238102
rect 331054 238046 331122 238102
rect 331178 238046 331248 238102
rect 330928 237978 331248 238046
rect 330928 237922 330998 237978
rect 331054 237922 331122 237978
rect 331178 237922 331248 237978
rect 330928 237888 331248 237922
rect 361648 238350 361968 238384
rect 361648 238294 361718 238350
rect 361774 238294 361842 238350
rect 361898 238294 361968 238350
rect 361648 238226 361968 238294
rect 361648 238170 361718 238226
rect 361774 238170 361842 238226
rect 361898 238170 361968 238226
rect 361648 238102 361968 238170
rect 361648 238046 361718 238102
rect 361774 238046 361842 238102
rect 361898 238046 361968 238102
rect 361648 237978 361968 238046
rect 361648 237922 361718 237978
rect 361774 237922 361842 237978
rect 361898 237922 361968 237978
rect 361648 237888 361968 237922
rect 392368 238350 392688 238384
rect 392368 238294 392438 238350
rect 392494 238294 392562 238350
rect 392618 238294 392688 238350
rect 392368 238226 392688 238294
rect 392368 238170 392438 238226
rect 392494 238170 392562 238226
rect 392618 238170 392688 238226
rect 392368 238102 392688 238170
rect 392368 238046 392438 238102
rect 392494 238046 392562 238102
rect 392618 238046 392688 238102
rect 392368 237978 392688 238046
rect 392368 237922 392438 237978
rect 392494 237922 392562 237978
rect 392618 237922 392688 237978
rect 392368 237888 392688 237922
rect 423088 238350 423408 238384
rect 423088 238294 423158 238350
rect 423214 238294 423282 238350
rect 423338 238294 423408 238350
rect 423088 238226 423408 238294
rect 423088 238170 423158 238226
rect 423214 238170 423282 238226
rect 423338 238170 423408 238226
rect 423088 238102 423408 238170
rect 423088 238046 423158 238102
rect 423214 238046 423282 238102
rect 423338 238046 423408 238102
rect 423088 237978 423408 238046
rect 423088 237922 423158 237978
rect 423214 237922 423282 237978
rect 423338 237922 423408 237978
rect 423088 237888 423408 237922
rect 453808 238350 454128 238384
rect 453808 238294 453878 238350
rect 453934 238294 454002 238350
rect 454058 238294 454128 238350
rect 453808 238226 454128 238294
rect 453808 238170 453878 238226
rect 453934 238170 454002 238226
rect 454058 238170 454128 238226
rect 453808 238102 454128 238170
rect 453808 238046 453878 238102
rect 453934 238046 454002 238102
rect 454058 238046 454128 238102
rect 453808 237978 454128 238046
rect 453808 237922 453878 237978
rect 453934 237922 454002 237978
rect 454058 237922 454128 237978
rect 453808 237888 454128 237922
rect 484528 238350 484848 238384
rect 484528 238294 484598 238350
rect 484654 238294 484722 238350
rect 484778 238294 484848 238350
rect 484528 238226 484848 238294
rect 484528 238170 484598 238226
rect 484654 238170 484722 238226
rect 484778 238170 484848 238226
rect 484528 238102 484848 238170
rect 484528 238046 484598 238102
rect 484654 238046 484722 238102
rect 484778 238046 484848 238102
rect 484528 237978 484848 238046
rect 484528 237922 484598 237978
rect 484654 237922 484722 237978
rect 484778 237922 484848 237978
rect 484528 237888 484848 237922
rect 515248 238350 515568 238384
rect 515248 238294 515318 238350
rect 515374 238294 515442 238350
rect 515498 238294 515568 238350
rect 515248 238226 515568 238294
rect 515248 238170 515318 238226
rect 515374 238170 515442 238226
rect 515498 238170 515568 238226
rect 515248 238102 515568 238170
rect 515248 238046 515318 238102
rect 515374 238046 515442 238102
rect 515498 238046 515568 238102
rect 515248 237978 515568 238046
rect 515248 237922 515318 237978
rect 515374 237922 515442 237978
rect 515498 237922 515568 237978
rect 515248 237888 515568 237922
rect 545968 238350 546288 238384
rect 545968 238294 546038 238350
rect 546094 238294 546162 238350
rect 546218 238294 546288 238350
rect 545968 238226 546288 238294
rect 545968 238170 546038 238226
rect 546094 238170 546162 238226
rect 546218 238170 546288 238226
rect 545968 238102 546288 238170
rect 545968 238046 546038 238102
rect 546094 238046 546162 238102
rect 546218 238046 546288 238102
rect 545968 237978 546288 238046
rect 545968 237922 546038 237978
rect 546094 237922 546162 237978
rect 546218 237922 546288 237978
rect 545968 237888 546288 237922
rect 561154 238350 561774 255922
rect 561154 238294 561250 238350
rect 561306 238294 561374 238350
rect 561430 238294 561498 238350
rect 561554 238294 561622 238350
rect 561678 238294 561774 238350
rect 561154 238226 561774 238294
rect 561154 238170 561250 238226
rect 561306 238170 561374 238226
rect 561430 238170 561498 238226
rect 561554 238170 561622 238226
rect 561678 238170 561774 238226
rect 561154 238102 561774 238170
rect 561154 238046 561250 238102
rect 561306 238046 561374 238102
rect 561430 238046 561498 238102
rect 561554 238046 561622 238102
rect 561678 238046 561774 238102
rect 561154 237978 561774 238046
rect 561154 237922 561250 237978
rect 561306 237922 561374 237978
rect 561430 237922 561498 237978
rect 561554 237922 561622 237978
rect 561678 237922 561774 237978
rect 131248 226350 131568 226384
rect 131248 226294 131318 226350
rect 131374 226294 131442 226350
rect 131498 226294 131568 226350
rect 131248 226226 131568 226294
rect 131248 226170 131318 226226
rect 131374 226170 131442 226226
rect 131498 226170 131568 226226
rect 131248 226102 131568 226170
rect 131248 226046 131318 226102
rect 131374 226046 131442 226102
rect 131498 226046 131568 226102
rect 131248 225978 131568 226046
rect 131248 225922 131318 225978
rect 131374 225922 131442 225978
rect 131498 225922 131568 225978
rect 131248 225888 131568 225922
rect 161968 226350 162288 226384
rect 161968 226294 162038 226350
rect 162094 226294 162162 226350
rect 162218 226294 162288 226350
rect 161968 226226 162288 226294
rect 161968 226170 162038 226226
rect 162094 226170 162162 226226
rect 162218 226170 162288 226226
rect 161968 226102 162288 226170
rect 161968 226046 162038 226102
rect 162094 226046 162162 226102
rect 162218 226046 162288 226102
rect 161968 225978 162288 226046
rect 161968 225922 162038 225978
rect 162094 225922 162162 225978
rect 162218 225922 162288 225978
rect 161968 225888 162288 225922
rect 192688 226350 193008 226384
rect 192688 226294 192758 226350
rect 192814 226294 192882 226350
rect 192938 226294 193008 226350
rect 192688 226226 193008 226294
rect 192688 226170 192758 226226
rect 192814 226170 192882 226226
rect 192938 226170 193008 226226
rect 192688 226102 193008 226170
rect 192688 226046 192758 226102
rect 192814 226046 192882 226102
rect 192938 226046 193008 226102
rect 192688 225978 193008 226046
rect 192688 225922 192758 225978
rect 192814 225922 192882 225978
rect 192938 225922 193008 225978
rect 192688 225888 193008 225922
rect 223408 226350 223728 226384
rect 223408 226294 223478 226350
rect 223534 226294 223602 226350
rect 223658 226294 223728 226350
rect 223408 226226 223728 226294
rect 223408 226170 223478 226226
rect 223534 226170 223602 226226
rect 223658 226170 223728 226226
rect 223408 226102 223728 226170
rect 223408 226046 223478 226102
rect 223534 226046 223602 226102
rect 223658 226046 223728 226102
rect 223408 225978 223728 226046
rect 223408 225922 223478 225978
rect 223534 225922 223602 225978
rect 223658 225922 223728 225978
rect 223408 225888 223728 225922
rect 254128 226350 254448 226384
rect 254128 226294 254198 226350
rect 254254 226294 254322 226350
rect 254378 226294 254448 226350
rect 254128 226226 254448 226294
rect 254128 226170 254198 226226
rect 254254 226170 254322 226226
rect 254378 226170 254448 226226
rect 254128 226102 254448 226170
rect 254128 226046 254198 226102
rect 254254 226046 254322 226102
rect 254378 226046 254448 226102
rect 254128 225978 254448 226046
rect 254128 225922 254198 225978
rect 254254 225922 254322 225978
rect 254378 225922 254448 225978
rect 254128 225888 254448 225922
rect 284848 226350 285168 226384
rect 284848 226294 284918 226350
rect 284974 226294 285042 226350
rect 285098 226294 285168 226350
rect 284848 226226 285168 226294
rect 284848 226170 284918 226226
rect 284974 226170 285042 226226
rect 285098 226170 285168 226226
rect 284848 226102 285168 226170
rect 284848 226046 284918 226102
rect 284974 226046 285042 226102
rect 285098 226046 285168 226102
rect 284848 225978 285168 226046
rect 284848 225922 284918 225978
rect 284974 225922 285042 225978
rect 285098 225922 285168 225978
rect 284848 225888 285168 225922
rect 315568 226350 315888 226384
rect 315568 226294 315638 226350
rect 315694 226294 315762 226350
rect 315818 226294 315888 226350
rect 315568 226226 315888 226294
rect 315568 226170 315638 226226
rect 315694 226170 315762 226226
rect 315818 226170 315888 226226
rect 315568 226102 315888 226170
rect 315568 226046 315638 226102
rect 315694 226046 315762 226102
rect 315818 226046 315888 226102
rect 315568 225978 315888 226046
rect 315568 225922 315638 225978
rect 315694 225922 315762 225978
rect 315818 225922 315888 225978
rect 315568 225888 315888 225922
rect 346288 226350 346608 226384
rect 346288 226294 346358 226350
rect 346414 226294 346482 226350
rect 346538 226294 346608 226350
rect 346288 226226 346608 226294
rect 346288 226170 346358 226226
rect 346414 226170 346482 226226
rect 346538 226170 346608 226226
rect 346288 226102 346608 226170
rect 346288 226046 346358 226102
rect 346414 226046 346482 226102
rect 346538 226046 346608 226102
rect 346288 225978 346608 226046
rect 346288 225922 346358 225978
rect 346414 225922 346482 225978
rect 346538 225922 346608 225978
rect 346288 225888 346608 225922
rect 377008 226350 377328 226384
rect 377008 226294 377078 226350
rect 377134 226294 377202 226350
rect 377258 226294 377328 226350
rect 377008 226226 377328 226294
rect 377008 226170 377078 226226
rect 377134 226170 377202 226226
rect 377258 226170 377328 226226
rect 377008 226102 377328 226170
rect 377008 226046 377078 226102
rect 377134 226046 377202 226102
rect 377258 226046 377328 226102
rect 377008 225978 377328 226046
rect 377008 225922 377078 225978
rect 377134 225922 377202 225978
rect 377258 225922 377328 225978
rect 377008 225888 377328 225922
rect 407728 226350 408048 226384
rect 407728 226294 407798 226350
rect 407854 226294 407922 226350
rect 407978 226294 408048 226350
rect 407728 226226 408048 226294
rect 407728 226170 407798 226226
rect 407854 226170 407922 226226
rect 407978 226170 408048 226226
rect 407728 226102 408048 226170
rect 407728 226046 407798 226102
rect 407854 226046 407922 226102
rect 407978 226046 408048 226102
rect 407728 225978 408048 226046
rect 407728 225922 407798 225978
rect 407854 225922 407922 225978
rect 407978 225922 408048 225978
rect 407728 225888 408048 225922
rect 438448 226350 438768 226384
rect 438448 226294 438518 226350
rect 438574 226294 438642 226350
rect 438698 226294 438768 226350
rect 438448 226226 438768 226294
rect 438448 226170 438518 226226
rect 438574 226170 438642 226226
rect 438698 226170 438768 226226
rect 438448 226102 438768 226170
rect 438448 226046 438518 226102
rect 438574 226046 438642 226102
rect 438698 226046 438768 226102
rect 438448 225978 438768 226046
rect 438448 225922 438518 225978
rect 438574 225922 438642 225978
rect 438698 225922 438768 225978
rect 438448 225888 438768 225922
rect 469168 226350 469488 226384
rect 469168 226294 469238 226350
rect 469294 226294 469362 226350
rect 469418 226294 469488 226350
rect 469168 226226 469488 226294
rect 469168 226170 469238 226226
rect 469294 226170 469362 226226
rect 469418 226170 469488 226226
rect 469168 226102 469488 226170
rect 469168 226046 469238 226102
rect 469294 226046 469362 226102
rect 469418 226046 469488 226102
rect 469168 225978 469488 226046
rect 469168 225922 469238 225978
rect 469294 225922 469362 225978
rect 469418 225922 469488 225978
rect 469168 225888 469488 225922
rect 499888 226350 500208 226384
rect 499888 226294 499958 226350
rect 500014 226294 500082 226350
rect 500138 226294 500208 226350
rect 499888 226226 500208 226294
rect 499888 226170 499958 226226
rect 500014 226170 500082 226226
rect 500138 226170 500208 226226
rect 499888 226102 500208 226170
rect 499888 226046 499958 226102
rect 500014 226046 500082 226102
rect 500138 226046 500208 226102
rect 499888 225978 500208 226046
rect 499888 225922 499958 225978
rect 500014 225922 500082 225978
rect 500138 225922 500208 225978
rect 499888 225888 500208 225922
rect 530608 226350 530928 226384
rect 530608 226294 530678 226350
rect 530734 226294 530802 226350
rect 530858 226294 530928 226350
rect 530608 226226 530928 226294
rect 530608 226170 530678 226226
rect 530734 226170 530802 226226
rect 530858 226170 530928 226226
rect 530608 226102 530928 226170
rect 530608 226046 530678 226102
rect 530734 226046 530802 226102
rect 530858 226046 530928 226102
rect 530608 225978 530928 226046
rect 530608 225922 530678 225978
rect 530734 225922 530802 225978
rect 530858 225922 530928 225978
rect 530608 225888 530928 225922
rect 111154 220294 111250 220350
rect 111306 220294 111374 220350
rect 111430 220294 111498 220350
rect 111554 220294 111622 220350
rect 111678 220294 111774 220350
rect 111154 220226 111774 220294
rect 111154 220170 111250 220226
rect 111306 220170 111374 220226
rect 111430 220170 111498 220226
rect 111554 220170 111622 220226
rect 111678 220170 111774 220226
rect 111154 220102 111774 220170
rect 111154 220046 111250 220102
rect 111306 220046 111374 220102
rect 111430 220046 111498 220102
rect 111554 220046 111622 220102
rect 111678 220046 111774 220102
rect 111154 219978 111774 220046
rect 111154 219922 111250 219978
rect 111306 219922 111374 219978
rect 111430 219922 111498 219978
rect 111554 219922 111622 219978
rect 111678 219922 111774 219978
rect 96874 208294 96970 208350
rect 97026 208294 97094 208350
rect 97150 208294 97218 208350
rect 97274 208294 97342 208350
rect 97398 208294 97494 208350
rect 96874 208226 97494 208294
rect 96874 208170 96970 208226
rect 97026 208170 97094 208226
rect 97150 208170 97218 208226
rect 97274 208170 97342 208226
rect 97398 208170 97494 208226
rect 96874 208102 97494 208170
rect 96874 208046 96970 208102
rect 97026 208046 97094 208102
rect 97150 208046 97218 208102
rect 97274 208046 97342 208102
rect 97398 208046 97494 208102
rect 96874 207978 97494 208046
rect 96874 207922 96970 207978
rect 97026 207922 97094 207978
rect 97150 207922 97218 207978
rect 97274 207922 97342 207978
rect 97398 207922 97494 207978
rect 96874 190350 97494 207922
rect 100528 208350 100848 208384
rect 100528 208294 100598 208350
rect 100654 208294 100722 208350
rect 100778 208294 100848 208350
rect 100528 208226 100848 208294
rect 100528 208170 100598 208226
rect 100654 208170 100722 208226
rect 100778 208170 100848 208226
rect 100528 208102 100848 208170
rect 100528 208046 100598 208102
rect 100654 208046 100722 208102
rect 100778 208046 100848 208102
rect 100528 207978 100848 208046
rect 100528 207922 100598 207978
rect 100654 207922 100722 207978
rect 100778 207922 100848 207978
rect 100528 207888 100848 207922
rect 111154 202350 111774 219922
rect 115888 220350 116208 220384
rect 115888 220294 115958 220350
rect 116014 220294 116082 220350
rect 116138 220294 116208 220350
rect 115888 220226 116208 220294
rect 115888 220170 115958 220226
rect 116014 220170 116082 220226
rect 116138 220170 116208 220226
rect 115888 220102 116208 220170
rect 115888 220046 115958 220102
rect 116014 220046 116082 220102
rect 116138 220046 116208 220102
rect 115888 219978 116208 220046
rect 115888 219922 115958 219978
rect 116014 219922 116082 219978
rect 116138 219922 116208 219978
rect 115888 219888 116208 219922
rect 146608 220350 146928 220384
rect 146608 220294 146678 220350
rect 146734 220294 146802 220350
rect 146858 220294 146928 220350
rect 146608 220226 146928 220294
rect 146608 220170 146678 220226
rect 146734 220170 146802 220226
rect 146858 220170 146928 220226
rect 146608 220102 146928 220170
rect 146608 220046 146678 220102
rect 146734 220046 146802 220102
rect 146858 220046 146928 220102
rect 146608 219978 146928 220046
rect 146608 219922 146678 219978
rect 146734 219922 146802 219978
rect 146858 219922 146928 219978
rect 146608 219888 146928 219922
rect 177328 220350 177648 220384
rect 177328 220294 177398 220350
rect 177454 220294 177522 220350
rect 177578 220294 177648 220350
rect 177328 220226 177648 220294
rect 177328 220170 177398 220226
rect 177454 220170 177522 220226
rect 177578 220170 177648 220226
rect 177328 220102 177648 220170
rect 177328 220046 177398 220102
rect 177454 220046 177522 220102
rect 177578 220046 177648 220102
rect 177328 219978 177648 220046
rect 177328 219922 177398 219978
rect 177454 219922 177522 219978
rect 177578 219922 177648 219978
rect 177328 219888 177648 219922
rect 208048 220350 208368 220384
rect 208048 220294 208118 220350
rect 208174 220294 208242 220350
rect 208298 220294 208368 220350
rect 208048 220226 208368 220294
rect 208048 220170 208118 220226
rect 208174 220170 208242 220226
rect 208298 220170 208368 220226
rect 208048 220102 208368 220170
rect 208048 220046 208118 220102
rect 208174 220046 208242 220102
rect 208298 220046 208368 220102
rect 208048 219978 208368 220046
rect 208048 219922 208118 219978
rect 208174 219922 208242 219978
rect 208298 219922 208368 219978
rect 208048 219888 208368 219922
rect 238768 220350 239088 220384
rect 238768 220294 238838 220350
rect 238894 220294 238962 220350
rect 239018 220294 239088 220350
rect 238768 220226 239088 220294
rect 238768 220170 238838 220226
rect 238894 220170 238962 220226
rect 239018 220170 239088 220226
rect 238768 220102 239088 220170
rect 238768 220046 238838 220102
rect 238894 220046 238962 220102
rect 239018 220046 239088 220102
rect 238768 219978 239088 220046
rect 238768 219922 238838 219978
rect 238894 219922 238962 219978
rect 239018 219922 239088 219978
rect 238768 219888 239088 219922
rect 269488 220350 269808 220384
rect 269488 220294 269558 220350
rect 269614 220294 269682 220350
rect 269738 220294 269808 220350
rect 269488 220226 269808 220294
rect 269488 220170 269558 220226
rect 269614 220170 269682 220226
rect 269738 220170 269808 220226
rect 269488 220102 269808 220170
rect 269488 220046 269558 220102
rect 269614 220046 269682 220102
rect 269738 220046 269808 220102
rect 269488 219978 269808 220046
rect 269488 219922 269558 219978
rect 269614 219922 269682 219978
rect 269738 219922 269808 219978
rect 269488 219888 269808 219922
rect 300208 220350 300528 220384
rect 300208 220294 300278 220350
rect 300334 220294 300402 220350
rect 300458 220294 300528 220350
rect 300208 220226 300528 220294
rect 300208 220170 300278 220226
rect 300334 220170 300402 220226
rect 300458 220170 300528 220226
rect 300208 220102 300528 220170
rect 300208 220046 300278 220102
rect 300334 220046 300402 220102
rect 300458 220046 300528 220102
rect 300208 219978 300528 220046
rect 300208 219922 300278 219978
rect 300334 219922 300402 219978
rect 300458 219922 300528 219978
rect 300208 219888 300528 219922
rect 330928 220350 331248 220384
rect 330928 220294 330998 220350
rect 331054 220294 331122 220350
rect 331178 220294 331248 220350
rect 330928 220226 331248 220294
rect 330928 220170 330998 220226
rect 331054 220170 331122 220226
rect 331178 220170 331248 220226
rect 330928 220102 331248 220170
rect 330928 220046 330998 220102
rect 331054 220046 331122 220102
rect 331178 220046 331248 220102
rect 330928 219978 331248 220046
rect 330928 219922 330998 219978
rect 331054 219922 331122 219978
rect 331178 219922 331248 219978
rect 330928 219888 331248 219922
rect 361648 220350 361968 220384
rect 361648 220294 361718 220350
rect 361774 220294 361842 220350
rect 361898 220294 361968 220350
rect 361648 220226 361968 220294
rect 361648 220170 361718 220226
rect 361774 220170 361842 220226
rect 361898 220170 361968 220226
rect 361648 220102 361968 220170
rect 361648 220046 361718 220102
rect 361774 220046 361842 220102
rect 361898 220046 361968 220102
rect 361648 219978 361968 220046
rect 361648 219922 361718 219978
rect 361774 219922 361842 219978
rect 361898 219922 361968 219978
rect 361648 219888 361968 219922
rect 392368 220350 392688 220384
rect 392368 220294 392438 220350
rect 392494 220294 392562 220350
rect 392618 220294 392688 220350
rect 392368 220226 392688 220294
rect 392368 220170 392438 220226
rect 392494 220170 392562 220226
rect 392618 220170 392688 220226
rect 392368 220102 392688 220170
rect 392368 220046 392438 220102
rect 392494 220046 392562 220102
rect 392618 220046 392688 220102
rect 392368 219978 392688 220046
rect 392368 219922 392438 219978
rect 392494 219922 392562 219978
rect 392618 219922 392688 219978
rect 392368 219888 392688 219922
rect 423088 220350 423408 220384
rect 423088 220294 423158 220350
rect 423214 220294 423282 220350
rect 423338 220294 423408 220350
rect 423088 220226 423408 220294
rect 423088 220170 423158 220226
rect 423214 220170 423282 220226
rect 423338 220170 423408 220226
rect 423088 220102 423408 220170
rect 423088 220046 423158 220102
rect 423214 220046 423282 220102
rect 423338 220046 423408 220102
rect 423088 219978 423408 220046
rect 423088 219922 423158 219978
rect 423214 219922 423282 219978
rect 423338 219922 423408 219978
rect 423088 219888 423408 219922
rect 453808 220350 454128 220384
rect 453808 220294 453878 220350
rect 453934 220294 454002 220350
rect 454058 220294 454128 220350
rect 453808 220226 454128 220294
rect 453808 220170 453878 220226
rect 453934 220170 454002 220226
rect 454058 220170 454128 220226
rect 453808 220102 454128 220170
rect 453808 220046 453878 220102
rect 453934 220046 454002 220102
rect 454058 220046 454128 220102
rect 453808 219978 454128 220046
rect 453808 219922 453878 219978
rect 453934 219922 454002 219978
rect 454058 219922 454128 219978
rect 453808 219888 454128 219922
rect 484528 220350 484848 220384
rect 484528 220294 484598 220350
rect 484654 220294 484722 220350
rect 484778 220294 484848 220350
rect 484528 220226 484848 220294
rect 484528 220170 484598 220226
rect 484654 220170 484722 220226
rect 484778 220170 484848 220226
rect 484528 220102 484848 220170
rect 484528 220046 484598 220102
rect 484654 220046 484722 220102
rect 484778 220046 484848 220102
rect 484528 219978 484848 220046
rect 484528 219922 484598 219978
rect 484654 219922 484722 219978
rect 484778 219922 484848 219978
rect 484528 219888 484848 219922
rect 515248 220350 515568 220384
rect 515248 220294 515318 220350
rect 515374 220294 515442 220350
rect 515498 220294 515568 220350
rect 515248 220226 515568 220294
rect 515248 220170 515318 220226
rect 515374 220170 515442 220226
rect 515498 220170 515568 220226
rect 515248 220102 515568 220170
rect 515248 220046 515318 220102
rect 515374 220046 515442 220102
rect 515498 220046 515568 220102
rect 515248 219978 515568 220046
rect 515248 219922 515318 219978
rect 515374 219922 515442 219978
rect 515498 219922 515568 219978
rect 515248 219888 515568 219922
rect 545968 220350 546288 220384
rect 545968 220294 546038 220350
rect 546094 220294 546162 220350
rect 546218 220294 546288 220350
rect 545968 220226 546288 220294
rect 545968 220170 546038 220226
rect 546094 220170 546162 220226
rect 546218 220170 546288 220226
rect 545968 220102 546288 220170
rect 545968 220046 546038 220102
rect 546094 220046 546162 220102
rect 546218 220046 546288 220102
rect 545968 219978 546288 220046
rect 545968 219922 546038 219978
rect 546094 219922 546162 219978
rect 546218 219922 546288 219978
rect 545968 219888 546288 219922
rect 561154 220350 561774 237922
rect 561154 220294 561250 220350
rect 561306 220294 561374 220350
rect 561430 220294 561498 220350
rect 561554 220294 561622 220350
rect 561678 220294 561774 220350
rect 561154 220226 561774 220294
rect 561154 220170 561250 220226
rect 561306 220170 561374 220226
rect 561430 220170 561498 220226
rect 561554 220170 561622 220226
rect 561678 220170 561774 220226
rect 561154 220102 561774 220170
rect 561154 220046 561250 220102
rect 561306 220046 561374 220102
rect 561430 220046 561498 220102
rect 561554 220046 561622 220102
rect 561678 220046 561774 220102
rect 561154 219978 561774 220046
rect 561154 219922 561250 219978
rect 561306 219922 561374 219978
rect 561430 219922 561498 219978
rect 561554 219922 561622 219978
rect 561678 219922 561774 219978
rect 131248 208350 131568 208384
rect 131248 208294 131318 208350
rect 131374 208294 131442 208350
rect 131498 208294 131568 208350
rect 131248 208226 131568 208294
rect 131248 208170 131318 208226
rect 131374 208170 131442 208226
rect 131498 208170 131568 208226
rect 131248 208102 131568 208170
rect 131248 208046 131318 208102
rect 131374 208046 131442 208102
rect 131498 208046 131568 208102
rect 131248 207978 131568 208046
rect 131248 207922 131318 207978
rect 131374 207922 131442 207978
rect 131498 207922 131568 207978
rect 131248 207888 131568 207922
rect 161968 208350 162288 208384
rect 161968 208294 162038 208350
rect 162094 208294 162162 208350
rect 162218 208294 162288 208350
rect 161968 208226 162288 208294
rect 161968 208170 162038 208226
rect 162094 208170 162162 208226
rect 162218 208170 162288 208226
rect 161968 208102 162288 208170
rect 161968 208046 162038 208102
rect 162094 208046 162162 208102
rect 162218 208046 162288 208102
rect 161968 207978 162288 208046
rect 161968 207922 162038 207978
rect 162094 207922 162162 207978
rect 162218 207922 162288 207978
rect 161968 207888 162288 207922
rect 192688 208350 193008 208384
rect 192688 208294 192758 208350
rect 192814 208294 192882 208350
rect 192938 208294 193008 208350
rect 192688 208226 193008 208294
rect 192688 208170 192758 208226
rect 192814 208170 192882 208226
rect 192938 208170 193008 208226
rect 192688 208102 193008 208170
rect 192688 208046 192758 208102
rect 192814 208046 192882 208102
rect 192938 208046 193008 208102
rect 192688 207978 193008 208046
rect 192688 207922 192758 207978
rect 192814 207922 192882 207978
rect 192938 207922 193008 207978
rect 192688 207888 193008 207922
rect 223408 208350 223728 208384
rect 223408 208294 223478 208350
rect 223534 208294 223602 208350
rect 223658 208294 223728 208350
rect 223408 208226 223728 208294
rect 223408 208170 223478 208226
rect 223534 208170 223602 208226
rect 223658 208170 223728 208226
rect 223408 208102 223728 208170
rect 223408 208046 223478 208102
rect 223534 208046 223602 208102
rect 223658 208046 223728 208102
rect 223408 207978 223728 208046
rect 223408 207922 223478 207978
rect 223534 207922 223602 207978
rect 223658 207922 223728 207978
rect 223408 207888 223728 207922
rect 254128 208350 254448 208384
rect 254128 208294 254198 208350
rect 254254 208294 254322 208350
rect 254378 208294 254448 208350
rect 254128 208226 254448 208294
rect 254128 208170 254198 208226
rect 254254 208170 254322 208226
rect 254378 208170 254448 208226
rect 254128 208102 254448 208170
rect 254128 208046 254198 208102
rect 254254 208046 254322 208102
rect 254378 208046 254448 208102
rect 254128 207978 254448 208046
rect 254128 207922 254198 207978
rect 254254 207922 254322 207978
rect 254378 207922 254448 207978
rect 254128 207888 254448 207922
rect 284848 208350 285168 208384
rect 284848 208294 284918 208350
rect 284974 208294 285042 208350
rect 285098 208294 285168 208350
rect 284848 208226 285168 208294
rect 284848 208170 284918 208226
rect 284974 208170 285042 208226
rect 285098 208170 285168 208226
rect 284848 208102 285168 208170
rect 284848 208046 284918 208102
rect 284974 208046 285042 208102
rect 285098 208046 285168 208102
rect 284848 207978 285168 208046
rect 284848 207922 284918 207978
rect 284974 207922 285042 207978
rect 285098 207922 285168 207978
rect 284848 207888 285168 207922
rect 315568 208350 315888 208384
rect 315568 208294 315638 208350
rect 315694 208294 315762 208350
rect 315818 208294 315888 208350
rect 315568 208226 315888 208294
rect 315568 208170 315638 208226
rect 315694 208170 315762 208226
rect 315818 208170 315888 208226
rect 315568 208102 315888 208170
rect 315568 208046 315638 208102
rect 315694 208046 315762 208102
rect 315818 208046 315888 208102
rect 315568 207978 315888 208046
rect 315568 207922 315638 207978
rect 315694 207922 315762 207978
rect 315818 207922 315888 207978
rect 315568 207888 315888 207922
rect 346288 208350 346608 208384
rect 346288 208294 346358 208350
rect 346414 208294 346482 208350
rect 346538 208294 346608 208350
rect 346288 208226 346608 208294
rect 346288 208170 346358 208226
rect 346414 208170 346482 208226
rect 346538 208170 346608 208226
rect 346288 208102 346608 208170
rect 346288 208046 346358 208102
rect 346414 208046 346482 208102
rect 346538 208046 346608 208102
rect 346288 207978 346608 208046
rect 346288 207922 346358 207978
rect 346414 207922 346482 207978
rect 346538 207922 346608 207978
rect 346288 207888 346608 207922
rect 377008 208350 377328 208384
rect 377008 208294 377078 208350
rect 377134 208294 377202 208350
rect 377258 208294 377328 208350
rect 377008 208226 377328 208294
rect 377008 208170 377078 208226
rect 377134 208170 377202 208226
rect 377258 208170 377328 208226
rect 377008 208102 377328 208170
rect 377008 208046 377078 208102
rect 377134 208046 377202 208102
rect 377258 208046 377328 208102
rect 377008 207978 377328 208046
rect 377008 207922 377078 207978
rect 377134 207922 377202 207978
rect 377258 207922 377328 207978
rect 377008 207888 377328 207922
rect 407728 208350 408048 208384
rect 407728 208294 407798 208350
rect 407854 208294 407922 208350
rect 407978 208294 408048 208350
rect 407728 208226 408048 208294
rect 407728 208170 407798 208226
rect 407854 208170 407922 208226
rect 407978 208170 408048 208226
rect 407728 208102 408048 208170
rect 407728 208046 407798 208102
rect 407854 208046 407922 208102
rect 407978 208046 408048 208102
rect 407728 207978 408048 208046
rect 407728 207922 407798 207978
rect 407854 207922 407922 207978
rect 407978 207922 408048 207978
rect 407728 207888 408048 207922
rect 438448 208350 438768 208384
rect 438448 208294 438518 208350
rect 438574 208294 438642 208350
rect 438698 208294 438768 208350
rect 438448 208226 438768 208294
rect 438448 208170 438518 208226
rect 438574 208170 438642 208226
rect 438698 208170 438768 208226
rect 438448 208102 438768 208170
rect 438448 208046 438518 208102
rect 438574 208046 438642 208102
rect 438698 208046 438768 208102
rect 438448 207978 438768 208046
rect 438448 207922 438518 207978
rect 438574 207922 438642 207978
rect 438698 207922 438768 207978
rect 438448 207888 438768 207922
rect 469168 208350 469488 208384
rect 469168 208294 469238 208350
rect 469294 208294 469362 208350
rect 469418 208294 469488 208350
rect 469168 208226 469488 208294
rect 469168 208170 469238 208226
rect 469294 208170 469362 208226
rect 469418 208170 469488 208226
rect 469168 208102 469488 208170
rect 469168 208046 469238 208102
rect 469294 208046 469362 208102
rect 469418 208046 469488 208102
rect 469168 207978 469488 208046
rect 469168 207922 469238 207978
rect 469294 207922 469362 207978
rect 469418 207922 469488 207978
rect 469168 207888 469488 207922
rect 499888 208350 500208 208384
rect 499888 208294 499958 208350
rect 500014 208294 500082 208350
rect 500138 208294 500208 208350
rect 499888 208226 500208 208294
rect 499888 208170 499958 208226
rect 500014 208170 500082 208226
rect 500138 208170 500208 208226
rect 499888 208102 500208 208170
rect 499888 208046 499958 208102
rect 500014 208046 500082 208102
rect 500138 208046 500208 208102
rect 499888 207978 500208 208046
rect 499888 207922 499958 207978
rect 500014 207922 500082 207978
rect 500138 207922 500208 207978
rect 499888 207888 500208 207922
rect 530608 208350 530928 208384
rect 530608 208294 530678 208350
rect 530734 208294 530802 208350
rect 530858 208294 530928 208350
rect 530608 208226 530928 208294
rect 530608 208170 530678 208226
rect 530734 208170 530802 208226
rect 530858 208170 530928 208226
rect 530608 208102 530928 208170
rect 530608 208046 530678 208102
rect 530734 208046 530802 208102
rect 530858 208046 530928 208102
rect 530608 207978 530928 208046
rect 530608 207922 530678 207978
rect 530734 207922 530802 207978
rect 530858 207922 530928 207978
rect 530608 207888 530928 207922
rect 111154 202294 111250 202350
rect 111306 202294 111374 202350
rect 111430 202294 111498 202350
rect 111554 202294 111622 202350
rect 111678 202294 111774 202350
rect 111154 202226 111774 202294
rect 111154 202170 111250 202226
rect 111306 202170 111374 202226
rect 111430 202170 111498 202226
rect 111554 202170 111622 202226
rect 111678 202170 111774 202226
rect 111154 202102 111774 202170
rect 111154 202046 111250 202102
rect 111306 202046 111374 202102
rect 111430 202046 111498 202102
rect 111554 202046 111622 202102
rect 111678 202046 111774 202102
rect 111154 201978 111774 202046
rect 111154 201922 111250 201978
rect 111306 201922 111374 201978
rect 111430 201922 111498 201978
rect 111554 201922 111622 201978
rect 111678 201922 111774 201978
rect 96874 190294 96970 190350
rect 97026 190294 97094 190350
rect 97150 190294 97218 190350
rect 97274 190294 97342 190350
rect 97398 190294 97494 190350
rect 96874 190226 97494 190294
rect 96874 190170 96970 190226
rect 97026 190170 97094 190226
rect 97150 190170 97218 190226
rect 97274 190170 97342 190226
rect 97398 190170 97494 190226
rect 96874 190102 97494 190170
rect 96874 190046 96970 190102
rect 97026 190046 97094 190102
rect 97150 190046 97218 190102
rect 97274 190046 97342 190102
rect 97398 190046 97494 190102
rect 96874 189978 97494 190046
rect 96874 189922 96970 189978
rect 97026 189922 97094 189978
rect 97150 189922 97218 189978
rect 97274 189922 97342 189978
rect 97398 189922 97494 189978
rect 96874 172350 97494 189922
rect 100528 190350 100848 190384
rect 100528 190294 100598 190350
rect 100654 190294 100722 190350
rect 100778 190294 100848 190350
rect 100528 190226 100848 190294
rect 100528 190170 100598 190226
rect 100654 190170 100722 190226
rect 100778 190170 100848 190226
rect 100528 190102 100848 190170
rect 100528 190046 100598 190102
rect 100654 190046 100722 190102
rect 100778 190046 100848 190102
rect 100528 189978 100848 190046
rect 100528 189922 100598 189978
rect 100654 189922 100722 189978
rect 100778 189922 100848 189978
rect 100528 189888 100848 189922
rect 111154 184350 111774 201922
rect 115888 202350 116208 202384
rect 115888 202294 115958 202350
rect 116014 202294 116082 202350
rect 116138 202294 116208 202350
rect 115888 202226 116208 202294
rect 115888 202170 115958 202226
rect 116014 202170 116082 202226
rect 116138 202170 116208 202226
rect 115888 202102 116208 202170
rect 115888 202046 115958 202102
rect 116014 202046 116082 202102
rect 116138 202046 116208 202102
rect 115888 201978 116208 202046
rect 115888 201922 115958 201978
rect 116014 201922 116082 201978
rect 116138 201922 116208 201978
rect 115888 201888 116208 201922
rect 146608 202350 146928 202384
rect 146608 202294 146678 202350
rect 146734 202294 146802 202350
rect 146858 202294 146928 202350
rect 146608 202226 146928 202294
rect 146608 202170 146678 202226
rect 146734 202170 146802 202226
rect 146858 202170 146928 202226
rect 146608 202102 146928 202170
rect 146608 202046 146678 202102
rect 146734 202046 146802 202102
rect 146858 202046 146928 202102
rect 146608 201978 146928 202046
rect 146608 201922 146678 201978
rect 146734 201922 146802 201978
rect 146858 201922 146928 201978
rect 146608 201888 146928 201922
rect 177328 202350 177648 202384
rect 177328 202294 177398 202350
rect 177454 202294 177522 202350
rect 177578 202294 177648 202350
rect 177328 202226 177648 202294
rect 177328 202170 177398 202226
rect 177454 202170 177522 202226
rect 177578 202170 177648 202226
rect 177328 202102 177648 202170
rect 177328 202046 177398 202102
rect 177454 202046 177522 202102
rect 177578 202046 177648 202102
rect 177328 201978 177648 202046
rect 177328 201922 177398 201978
rect 177454 201922 177522 201978
rect 177578 201922 177648 201978
rect 177328 201888 177648 201922
rect 208048 202350 208368 202384
rect 208048 202294 208118 202350
rect 208174 202294 208242 202350
rect 208298 202294 208368 202350
rect 208048 202226 208368 202294
rect 208048 202170 208118 202226
rect 208174 202170 208242 202226
rect 208298 202170 208368 202226
rect 208048 202102 208368 202170
rect 208048 202046 208118 202102
rect 208174 202046 208242 202102
rect 208298 202046 208368 202102
rect 208048 201978 208368 202046
rect 208048 201922 208118 201978
rect 208174 201922 208242 201978
rect 208298 201922 208368 201978
rect 208048 201888 208368 201922
rect 238768 202350 239088 202384
rect 238768 202294 238838 202350
rect 238894 202294 238962 202350
rect 239018 202294 239088 202350
rect 238768 202226 239088 202294
rect 238768 202170 238838 202226
rect 238894 202170 238962 202226
rect 239018 202170 239088 202226
rect 238768 202102 239088 202170
rect 238768 202046 238838 202102
rect 238894 202046 238962 202102
rect 239018 202046 239088 202102
rect 238768 201978 239088 202046
rect 238768 201922 238838 201978
rect 238894 201922 238962 201978
rect 239018 201922 239088 201978
rect 238768 201888 239088 201922
rect 269488 202350 269808 202384
rect 269488 202294 269558 202350
rect 269614 202294 269682 202350
rect 269738 202294 269808 202350
rect 269488 202226 269808 202294
rect 269488 202170 269558 202226
rect 269614 202170 269682 202226
rect 269738 202170 269808 202226
rect 269488 202102 269808 202170
rect 269488 202046 269558 202102
rect 269614 202046 269682 202102
rect 269738 202046 269808 202102
rect 269488 201978 269808 202046
rect 269488 201922 269558 201978
rect 269614 201922 269682 201978
rect 269738 201922 269808 201978
rect 269488 201888 269808 201922
rect 300208 202350 300528 202384
rect 300208 202294 300278 202350
rect 300334 202294 300402 202350
rect 300458 202294 300528 202350
rect 300208 202226 300528 202294
rect 300208 202170 300278 202226
rect 300334 202170 300402 202226
rect 300458 202170 300528 202226
rect 300208 202102 300528 202170
rect 300208 202046 300278 202102
rect 300334 202046 300402 202102
rect 300458 202046 300528 202102
rect 300208 201978 300528 202046
rect 300208 201922 300278 201978
rect 300334 201922 300402 201978
rect 300458 201922 300528 201978
rect 300208 201888 300528 201922
rect 330928 202350 331248 202384
rect 330928 202294 330998 202350
rect 331054 202294 331122 202350
rect 331178 202294 331248 202350
rect 330928 202226 331248 202294
rect 330928 202170 330998 202226
rect 331054 202170 331122 202226
rect 331178 202170 331248 202226
rect 330928 202102 331248 202170
rect 330928 202046 330998 202102
rect 331054 202046 331122 202102
rect 331178 202046 331248 202102
rect 330928 201978 331248 202046
rect 330928 201922 330998 201978
rect 331054 201922 331122 201978
rect 331178 201922 331248 201978
rect 330928 201888 331248 201922
rect 361648 202350 361968 202384
rect 361648 202294 361718 202350
rect 361774 202294 361842 202350
rect 361898 202294 361968 202350
rect 361648 202226 361968 202294
rect 361648 202170 361718 202226
rect 361774 202170 361842 202226
rect 361898 202170 361968 202226
rect 361648 202102 361968 202170
rect 361648 202046 361718 202102
rect 361774 202046 361842 202102
rect 361898 202046 361968 202102
rect 361648 201978 361968 202046
rect 361648 201922 361718 201978
rect 361774 201922 361842 201978
rect 361898 201922 361968 201978
rect 361648 201888 361968 201922
rect 392368 202350 392688 202384
rect 392368 202294 392438 202350
rect 392494 202294 392562 202350
rect 392618 202294 392688 202350
rect 392368 202226 392688 202294
rect 392368 202170 392438 202226
rect 392494 202170 392562 202226
rect 392618 202170 392688 202226
rect 392368 202102 392688 202170
rect 392368 202046 392438 202102
rect 392494 202046 392562 202102
rect 392618 202046 392688 202102
rect 392368 201978 392688 202046
rect 392368 201922 392438 201978
rect 392494 201922 392562 201978
rect 392618 201922 392688 201978
rect 392368 201888 392688 201922
rect 423088 202350 423408 202384
rect 423088 202294 423158 202350
rect 423214 202294 423282 202350
rect 423338 202294 423408 202350
rect 423088 202226 423408 202294
rect 423088 202170 423158 202226
rect 423214 202170 423282 202226
rect 423338 202170 423408 202226
rect 423088 202102 423408 202170
rect 423088 202046 423158 202102
rect 423214 202046 423282 202102
rect 423338 202046 423408 202102
rect 423088 201978 423408 202046
rect 423088 201922 423158 201978
rect 423214 201922 423282 201978
rect 423338 201922 423408 201978
rect 423088 201888 423408 201922
rect 453808 202350 454128 202384
rect 453808 202294 453878 202350
rect 453934 202294 454002 202350
rect 454058 202294 454128 202350
rect 453808 202226 454128 202294
rect 453808 202170 453878 202226
rect 453934 202170 454002 202226
rect 454058 202170 454128 202226
rect 453808 202102 454128 202170
rect 453808 202046 453878 202102
rect 453934 202046 454002 202102
rect 454058 202046 454128 202102
rect 453808 201978 454128 202046
rect 453808 201922 453878 201978
rect 453934 201922 454002 201978
rect 454058 201922 454128 201978
rect 453808 201888 454128 201922
rect 484528 202350 484848 202384
rect 484528 202294 484598 202350
rect 484654 202294 484722 202350
rect 484778 202294 484848 202350
rect 484528 202226 484848 202294
rect 484528 202170 484598 202226
rect 484654 202170 484722 202226
rect 484778 202170 484848 202226
rect 484528 202102 484848 202170
rect 484528 202046 484598 202102
rect 484654 202046 484722 202102
rect 484778 202046 484848 202102
rect 484528 201978 484848 202046
rect 484528 201922 484598 201978
rect 484654 201922 484722 201978
rect 484778 201922 484848 201978
rect 484528 201888 484848 201922
rect 515248 202350 515568 202384
rect 515248 202294 515318 202350
rect 515374 202294 515442 202350
rect 515498 202294 515568 202350
rect 515248 202226 515568 202294
rect 515248 202170 515318 202226
rect 515374 202170 515442 202226
rect 515498 202170 515568 202226
rect 515248 202102 515568 202170
rect 515248 202046 515318 202102
rect 515374 202046 515442 202102
rect 515498 202046 515568 202102
rect 515248 201978 515568 202046
rect 515248 201922 515318 201978
rect 515374 201922 515442 201978
rect 515498 201922 515568 201978
rect 515248 201888 515568 201922
rect 545968 202350 546288 202384
rect 545968 202294 546038 202350
rect 546094 202294 546162 202350
rect 546218 202294 546288 202350
rect 545968 202226 546288 202294
rect 545968 202170 546038 202226
rect 546094 202170 546162 202226
rect 546218 202170 546288 202226
rect 545968 202102 546288 202170
rect 545968 202046 546038 202102
rect 546094 202046 546162 202102
rect 546218 202046 546288 202102
rect 545968 201978 546288 202046
rect 545968 201922 546038 201978
rect 546094 201922 546162 201978
rect 546218 201922 546288 201978
rect 545968 201888 546288 201922
rect 561154 202350 561774 219922
rect 561154 202294 561250 202350
rect 561306 202294 561374 202350
rect 561430 202294 561498 202350
rect 561554 202294 561622 202350
rect 561678 202294 561774 202350
rect 561154 202226 561774 202294
rect 561154 202170 561250 202226
rect 561306 202170 561374 202226
rect 561430 202170 561498 202226
rect 561554 202170 561622 202226
rect 561678 202170 561774 202226
rect 561154 202102 561774 202170
rect 561154 202046 561250 202102
rect 561306 202046 561374 202102
rect 561430 202046 561498 202102
rect 561554 202046 561622 202102
rect 561678 202046 561774 202102
rect 561154 201978 561774 202046
rect 561154 201922 561250 201978
rect 561306 201922 561374 201978
rect 561430 201922 561498 201978
rect 561554 201922 561622 201978
rect 561678 201922 561774 201978
rect 131248 190350 131568 190384
rect 131248 190294 131318 190350
rect 131374 190294 131442 190350
rect 131498 190294 131568 190350
rect 131248 190226 131568 190294
rect 131248 190170 131318 190226
rect 131374 190170 131442 190226
rect 131498 190170 131568 190226
rect 131248 190102 131568 190170
rect 131248 190046 131318 190102
rect 131374 190046 131442 190102
rect 131498 190046 131568 190102
rect 131248 189978 131568 190046
rect 131248 189922 131318 189978
rect 131374 189922 131442 189978
rect 131498 189922 131568 189978
rect 131248 189888 131568 189922
rect 161968 190350 162288 190384
rect 161968 190294 162038 190350
rect 162094 190294 162162 190350
rect 162218 190294 162288 190350
rect 161968 190226 162288 190294
rect 161968 190170 162038 190226
rect 162094 190170 162162 190226
rect 162218 190170 162288 190226
rect 161968 190102 162288 190170
rect 161968 190046 162038 190102
rect 162094 190046 162162 190102
rect 162218 190046 162288 190102
rect 161968 189978 162288 190046
rect 161968 189922 162038 189978
rect 162094 189922 162162 189978
rect 162218 189922 162288 189978
rect 161968 189888 162288 189922
rect 192688 190350 193008 190384
rect 192688 190294 192758 190350
rect 192814 190294 192882 190350
rect 192938 190294 193008 190350
rect 192688 190226 193008 190294
rect 192688 190170 192758 190226
rect 192814 190170 192882 190226
rect 192938 190170 193008 190226
rect 192688 190102 193008 190170
rect 192688 190046 192758 190102
rect 192814 190046 192882 190102
rect 192938 190046 193008 190102
rect 192688 189978 193008 190046
rect 192688 189922 192758 189978
rect 192814 189922 192882 189978
rect 192938 189922 193008 189978
rect 192688 189888 193008 189922
rect 223408 190350 223728 190384
rect 223408 190294 223478 190350
rect 223534 190294 223602 190350
rect 223658 190294 223728 190350
rect 223408 190226 223728 190294
rect 223408 190170 223478 190226
rect 223534 190170 223602 190226
rect 223658 190170 223728 190226
rect 223408 190102 223728 190170
rect 223408 190046 223478 190102
rect 223534 190046 223602 190102
rect 223658 190046 223728 190102
rect 223408 189978 223728 190046
rect 223408 189922 223478 189978
rect 223534 189922 223602 189978
rect 223658 189922 223728 189978
rect 223408 189888 223728 189922
rect 254128 190350 254448 190384
rect 254128 190294 254198 190350
rect 254254 190294 254322 190350
rect 254378 190294 254448 190350
rect 254128 190226 254448 190294
rect 254128 190170 254198 190226
rect 254254 190170 254322 190226
rect 254378 190170 254448 190226
rect 254128 190102 254448 190170
rect 254128 190046 254198 190102
rect 254254 190046 254322 190102
rect 254378 190046 254448 190102
rect 254128 189978 254448 190046
rect 254128 189922 254198 189978
rect 254254 189922 254322 189978
rect 254378 189922 254448 189978
rect 254128 189888 254448 189922
rect 284848 190350 285168 190384
rect 284848 190294 284918 190350
rect 284974 190294 285042 190350
rect 285098 190294 285168 190350
rect 284848 190226 285168 190294
rect 284848 190170 284918 190226
rect 284974 190170 285042 190226
rect 285098 190170 285168 190226
rect 284848 190102 285168 190170
rect 284848 190046 284918 190102
rect 284974 190046 285042 190102
rect 285098 190046 285168 190102
rect 284848 189978 285168 190046
rect 284848 189922 284918 189978
rect 284974 189922 285042 189978
rect 285098 189922 285168 189978
rect 284848 189888 285168 189922
rect 315568 190350 315888 190384
rect 315568 190294 315638 190350
rect 315694 190294 315762 190350
rect 315818 190294 315888 190350
rect 315568 190226 315888 190294
rect 315568 190170 315638 190226
rect 315694 190170 315762 190226
rect 315818 190170 315888 190226
rect 315568 190102 315888 190170
rect 315568 190046 315638 190102
rect 315694 190046 315762 190102
rect 315818 190046 315888 190102
rect 315568 189978 315888 190046
rect 315568 189922 315638 189978
rect 315694 189922 315762 189978
rect 315818 189922 315888 189978
rect 315568 189888 315888 189922
rect 346288 190350 346608 190384
rect 346288 190294 346358 190350
rect 346414 190294 346482 190350
rect 346538 190294 346608 190350
rect 346288 190226 346608 190294
rect 346288 190170 346358 190226
rect 346414 190170 346482 190226
rect 346538 190170 346608 190226
rect 346288 190102 346608 190170
rect 346288 190046 346358 190102
rect 346414 190046 346482 190102
rect 346538 190046 346608 190102
rect 346288 189978 346608 190046
rect 346288 189922 346358 189978
rect 346414 189922 346482 189978
rect 346538 189922 346608 189978
rect 346288 189888 346608 189922
rect 377008 190350 377328 190384
rect 377008 190294 377078 190350
rect 377134 190294 377202 190350
rect 377258 190294 377328 190350
rect 377008 190226 377328 190294
rect 377008 190170 377078 190226
rect 377134 190170 377202 190226
rect 377258 190170 377328 190226
rect 377008 190102 377328 190170
rect 377008 190046 377078 190102
rect 377134 190046 377202 190102
rect 377258 190046 377328 190102
rect 377008 189978 377328 190046
rect 377008 189922 377078 189978
rect 377134 189922 377202 189978
rect 377258 189922 377328 189978
rect 377008 189888 377328 189922
rect 407728 190350 408048 190384
rect 407728 190294 407798 190350
rect 407854 190294 407922 190350
rect 407978 190294 408048 190350
rect 407728 190226 408048 190294
rect 407728 190170 407798 190226
rect 407854 190170 407922 190226
rect 407978 190170 408048 190226
rect 407728 190102 408048 190170
rect 407728 190046 407798 190102
rect 407854 190046 407922 190102
rect 407978 190046 408048 190102
rect 407728 189978 408048 190046
rect 407728 189922 407798 189978
rect 407854 189922 407922 189978
rect 407978 189922 408048 189978
rect 407728 189888 408048 189922
rect 438448 190350 438768 190384
rect 438448 190294 438518 190350
rect 438574 190294 438642 190350
rect 438698 190294 438768 190350
rect 438448 190226 438768 190294
rect 438448 190170 438518 190226
rect 438574 190170 438642 190226
rect 438698 190170 438768 190226
rect 438448 190102 438768 190170
rect 438448 190046 438518 190102
rect 438574 190046 438642 190102
rect 438698 190046 438768 190102
rect 438448 189978 438768 190046
rect 438448 189922 438518 189978
rect 438574 189922 438642 189978
rect 438698 189922 438768 189978
rect 438448 189888 438768 189922
rect 469168 190350 469488 190384
rect 469168 190294 469238 190350
rect 469294 190294 469362 190350
rect 469418 190294 469488 190350
rect 469168 190226 469488 190294
rect 469168 190170 469238 190226
rect 469294 190170 469362 190226
rect 469418 190170 469488 190226
rect 469168 190102 469488 190170
rect 469168 190046 469238 190102
rect 469294 190046 469362 190102
rect 469418 190046 469488 190102
rect 469168 189978 469488 190046
rect 469168 189922 469238 189978
rect 469294 189922 469362 189978
rect 469418 189922 469488 189978
rect 469168 189888 469488 189922
rect 499888 190350 500208 190384
rect 499888 190294 499958 190350
rect 500014 190294 500082 190350
rect 500138 190294 500208 190350
rect 499888 190226 500208 190294
rect 499888 190170 499958 190226
rect 500014 190170 500082 190226
rect 500138 190170 500208 190226
rect 499888 190102 500208 190170
rect 499888 190046 499958 190102
rect 500014 190046 500082 190102
rect 500138 190046 500208 190102
rect 499888 189978 500208 190046
rect 499888 189922 499958 189978
rect 500014 189922 500082 189978
rect 500138 189922 500208 189978
rect 499888 189888 500208 189922
rect 530608 190350 530928 190384
rect 530608 190294 530678 190350
rect 530734 190294 530802 190350
rect 530858 190294 530928 190350
rect 530608 190226 530928 190294
rect 530608 190170 530678 190226
rect 530734 190170 530802 190226
rect 530858 190170 530928 190226
rect 530608 190102 530928 190170
rect 530608 190046 530678 190102
rect 530734 190046 530802 190102
rect 530858 190046 530928 190102
rect 530608 189978 530928 190046
rect 530608 189922 530678 189978
rect 530734 189922 530802 189978
rect 530858 189922 530928 189978
rect 530608 189888 530928 189922
rect 111154 184294 111250 184350
rect 111306 184294 111374 184350
rect 111430 184294 111498 184350
rect 111554 184294 111622 184350
rect 111678 184294 111774 184350
rect 111154 184226 111774 184294
rect 111154 184170 111250 184226
rect 111306 184170 111374 184226
rect 111430 184170 111498 184226
rect 111554 184170 111622 184226
rect 111678 184170 111774 184226
rect 111154 184102 111774 184170
rect 111154 184046 111250 184102
rect 111306 184046 111374 184102
rect 111430 184046 111498 184102
rect 111554 184046 111622 184102
rect 111678 184046 111774 184102
rect 111154 183978 111774 184046
rect 111154 183922 111250 183978
rect 111306 183922 111374 183978
rect 111430 183922 111498 183978
rect 111554 183922 111622 183978
rect 111678 183922 111774 183978
rect 96874 172294 96970 172350
rect 97026 172294 97094 172350
rect 97150 172294 97218 172350
rect 97274 172294 97342 172350
rect 97398 172294 97494 172350
rect 96874 172226 97494 172294
rect 96874 172170 96970 172226
rect 97026 172170 97094 172226
rect 97150 172170 97218 172226
rect 97274 172170 97342 172226
rect 97398 172170 97494 172226
rect 96874 172102 97494 172170
rect 96874 172046 96970 172102
rect 97026 172046 97094 172102
rect 97150 172046 97218 172102
rect 97274 172046 97342 172102
rect 97398 172046 97494 172102
rect 96874 171978 97494 172046
rect 96874 171922 96970 171978
rect 97026 171922 97094 171978
rect 97150 171922 97218 171978
rect 97274 171922 97342 171978
rect 97398 171922 97494 171978
rect 96874 154350 97494 171922
rect 100528 172350 100848 172384
rect 100528 172294 100598 172350
rect 100654 172294 100722 172350
rect 100778 172294 100848 172350
rect 100528 172226 100848 172294
rect 100528 172170 100598 172226
rect 100654 172170 100722 172226
rect 100778 172170 100848 172226
rect 100528 172102 100848 172170
rect 100528 172046 100598 172102
rect 100654 172046 100722 172102
rect 100778 172046 100848 172102
rect 100528 171978 100848 172046
rect 100528 171922 100598 171978
rect 100654 171922 100722 171978
rect 100778 171922 100848 171978
rect 100528 171888 100848 171922
rect 111154 166350 111774 183922
rect 115888 184350 116208 184384
rect 115888 184294 115958 184350
rect 116014 184294 116082 184350
rect 116138 184294 116208 184350
rect 115888 184226 116208 184294
rect 115888 184170 115958 184226
rect 116014 184170 116082 184226
rect 116138 184170 116208 184226
rect 115888 184102 116208 184170
rect 115888 184046 115958 184102
rect 116014 184046 116082 184102
rect 116138 184046 116208 184102
rect 115888 183978 116208 184046
rect 115888 183922 115958 183978
rect 116014 183922 116082 183978
rect 116138 183922 116208 183978
rect 115888 183888 116208 183922
rect 146608 184350 146928 184384
rect 146608 184294 146678 184350
rect 146734 184294 146802 184350
rect 146858 184294 146928 184350
rect 146608 184226 146928 184294
rect 146608 184170 146678 184226
rect 146734 184170 146802 184226
rect 146858 184170 146928 184226
rect 146608 184102 146928 184170
rect 146608 184046 146678 184102
rect 146734 184046 146802 184102
rect 146858 184046 146928 184102
rect 146608 183978 146928 184046
rect 146608 183922 146678 183978
rect 146734 183922 146802 183978
rect 146858 183922 146928 183978
rect 146608 183888 146928 183922
rect 177328 184350 177648 184384
rect 177328 184294 177398 184350
rect 177454 184294 177522 184350
rect 177578 184294 177648 184350
rect 177328 184226 177648 184294
rect 177328 184170 177398 184226
rect 177454 184170 177522 184226
rect 177578 184170 177648 184226
rect 177328 184102 177648 184170
rect 177328 184046 177398 184102
rect 177454 184046 177522 184102
rect 177578 184046 177648 184102
rect 177328 183978 177648 184046
rect 177328 183922 177398 183978
rect 177454 183922 177522 183978
rect 177578 183922 177648 183978
rect 177328 183888 177648 183922
rect 208048 184350 208368 184384
rect 208048 184294 208118 184350
rect 208174 184294 208242 184350
rect 208298 184294 208368 184350
rect 208048 184226 208368 184294
rect 208048 184170 208118 184226
rect 208174 184170 208242 184226
rect 208298 184170 208368 184226
rect 208048 184102 208368 184170
rect 208048 184046 208118 184102
rect 208174 184046 208242 184102
rect 208298 184046 208368 184102
rect 208048 183978 208368 184046
rect 208048 183922 208118 183978
rect 208174 183922 208242 183978
rect 208298 183922 208368 183978
rect 208048 183888 208368 183922
rect 238768 184350 239088 184384
rect 238768 184294 238838 184350
rect 238894 184294 238962 184350
rect 239018 184294 239088 184350
rect 238768 184226 239088 184294
rect 238768 184170 238838 184226
rect 238894 184170 238962 184226
rect 239018 184170 239088 184226
rect 238768 184102 239088 184170
rect 238768 184046 238838 184102
rect 238894 184046 238962 184102
rect 239018 184046 239088 184102
rect 238768 183978 239088 184046
rect 238768 183922 238838 183978
rect 238894 183922 238962 183978
rect 239018 183922 239088 183978
rect 238768 183888 239088 183922
rect 269488 184350 269808 184384
rect 269488 184294 269558 184350
rect 269614 184294 269682 184350
rect 269738 184294 269808 184350
rect 269488 184226 269808 184294
rect 269488 184170 269558 184226
rect 269614 184170 269682 184226
rect 269738 184170 269808 184226
rect 269488 184102 269808 184170
rect 269488 184046 269558 184102
rect 269614 184046 269682 184102
rect 269738 184046 269808 184102
rect 269488 183978 269808 184046
rect 269488 183922 269558 183978
rect 269614 183922 269682 183978
rect 269738 183922 269808 183978
rect 269488 183888 269808 183922
rect 300208 184350 300528 184384
rect 300208 184294 300278 184350
rect 300334 184294 300402 184350
rect 300458 184294 300528 184350
rect 300208 184226 300528 184294
rect 300208 184170 300278 184226
rect 300334 184170 300402 184226
rect 300458 184170 300528 184226
rect 300208 184102 300528 184170
rect 300208 184046 300278 184102
rect 300334 184046 300402 184102
rect 300458 184046 300528 184102
rect 300208 183978 300528 184046
rect 300208 183922 300278 183978
rect 300334 183922 300402 183978
rect 300458 183922 300528 183978
rect 300208 183888 300528 183922
rect 330928 184350 331248 184384
rect 330928 184294 330998 184350
rect 331054 184294 331122 184350
rect 331178 184294 331248 184350
rect 330928 184226 331248 184294
rect 330928 184170 330998 184226
rect 331054 184170 331122 184226
rect 331178 184170 331248 184226
rect 330928 184102 331248 184170
rect 330928 184046 330998 184102
rect 331054 184046 331122 184102
rect 331178 184046 331248 184102
rect 330928 183978 331248 184046
rect 330928 183922 330998 183978
rect 331054 183922 331122 183978
rect 331178 183922 331248 183978
rect 330928 183888 331248 183922
rect 361648 184350 361968 184384
rect 361648 184294 361718 184350
rect 361774 184294 361842 184350
rect 361898 184294 361968 184350
rect 361648 184226 361968 184294
rect 361648 184170 361718 184226
rect 361774 184170 361842 184226
rect 361898 184170 361968 184226
rect 361648 184102 361968 184170
rect 361648 184046 361718 184102
rect 361774 184046 361842 184102
rect 361898 184046 361968 184102
rect 361648 183978 361968 184046
rect 361648 183922 361718 183978
rect 361774 183922 361842 183978
rect 361898 183922 361968 183978
rect 361648 183888 361968 183922
rect 392368 184350 392688 184384
rect 392368 184294 392438 184350
rect 392494 184294 392562 184350
rect 392618 184294 392688 184350
rect 392368 184226 392688 184294
rect 392368 184170 392438 184226
rect 392494 184170 392562 184226
rect 392618 184170 392688 184226
rect 392368 184102 392688 184170
rect 392368 184046 392438 184102
rect 392494 184046 392562 184102
rect 392618 184046 392688 184102
rect 392368 183978 392688 184046
rect 392368 183922 392438 183978
rect 392494 183922 392562 183978
rect 392618 183922 392688 183978
rect 392368 183888 392688 183922
rect 423088 184350 423408 184384
rect 423088 184294 423158 184350
rect 423214 184294 423282 184350
rect 423338 184294 423408 184350
rect 423088 184226 423408 184294
rect 423088 184170 423158 184226
rect 423214 184170 423282 184226
rect 423338 184170 423408 184226
rect 423088 184102 423408 184170
rect 423088 184046 423158 184102
rect 423214 184046 423282 184102
rect 423338 184046 423408 184102
rect 423088 183978 423408 184046
rect 423088 183922 423158 183978
rect 423214 183922 423282 183978
rect 423338 183922 423408 183978
rect 423088 183888 423408 183922
rect 453808 184350 454128 184384
rect 453808 184294 453878 184350
rect 453934 184294 454002 184350
rect 454058 184294 454128 184350
rect 453808 184226 454128 184294
rect 453808 184170 453878 184226
rect 453934 184170 454002 184226
rect 454058 184170 454128 184226
rect 453808 184102 454128 184170
rect 453808 184046 453878 184102
rect 453934 184046 454002 184102
rect 454058 184046 454128 184102
rect 453808 183978 454128 184046
rect 453808 183922 453878 183978
rect 453934 183922 454002 183978
rect 454058 183922 454128 183978
rect 453808 183888 454128 183922
rect 484528 184350 484848 184384
rect 484528 184294 484598 184350
rect 484654 184294 484722 184350
rect 484778 184294 484848 184350
rect 484528 184226 484848 184294
rect 484528 184170 484598 184226
rect 484654 184170 484722 184226
rect 484778 184170 484848 184226
rect 484528 184102 484848 184170
rect 484528 184046 484598 184102
rect 484654 184046 484722 184102
rect 484778 184046 484848 184102
rect 484528 183978 484848 184046
rect 484528 183922 484598 183978
rect 484654 183922 484722 183978
rect 484778 183922 484848 183978
rect 484528 183888 484848 183922
rect 515248 184350 515568 184384
rect 515248 184294 515318 184350
rect 515374 184294 515442 184350
rect 515498 184294 515568 184350
rect 515248 184226 515568 184294
rect 515248 184170 515318 184226
rect 515374 184170 515442 184226
rect 515498 184170 515568 184226
rect 515248 184102 515568 184170
rect 515248 184046 515318 184102
rect 515374 184046 515442 184102
rect 515498 184046 515568 184102
rect 515248 183978 515568 184046
rect 515248 183922 515318 183978
rect 515374 183922 515442 183978
rect 515498 183922 515568 183978
rect 515248 183888 515568 183922
rect 545968 184350 546288 184384
rect 545968 184294 546038 184350
rect 546094 184294 546162 184350
rect 546218 184294 546288 184350
rect 545968 184226 546288 184294
rect 545968 184170 546038 184226
rect 546094 184170 546162 184226
rect 546218 184170 546288 184226
rect 545968 184102 546288 184170
rect 545968 184046 546038 184102
rect 546094 184046 546162 184102
rect 546218 184046 546288 184102
rect 545968 183978 546288 184046
rect 545968 183922 546038 183978
rect 546094 183922 546162 183978
rect 546218 183922 546288 183978
rect 545968 183888 546288 183922
rect 561154 184350 561774 201922
rect 561154 184294 561250 184350
rect 561306 184294 561374 184350
rect 561430 184294 561498 184350
rect 561554 184294 561622 184350
rect 561678 184294 561774 184350
rect 561154 184226 561774 184294
rect 561154 184170 561250 184226
rect 561306 184170 561374 184226
rect 561430 184170 561498 184226
rect 561554 184170 561622 184226
rect 561678 184170 561774 184226
rect 561154 184102 561774 184170
rect 561154 184046 561250 184102
rect 561306 184046 561374 184102
rect 561430 184046 561498 184102
rect 561554 184046 561622 184102
rect 561678 184046 561774 184102
rect 561154 183978 561774 184046
rect 561154 183922 561250 183978
rect 561306 183922 561374 183978
rect 561430 183922 561498 183978
rect 561554 183922 561622 183978
rect 561678 183922 561774 183978
rect 131248 172350 131568 172384
rect 131248 172294 131318 172350
rect 131374 172294 131442 172350
rect 131498 172294 131568 172350
rect 131248 172226 131568 172294
rect 131248 172170 131318 172226
rect 131374 172170 131442 172226
rect 131498 172170 131568 172226
rect 131248 172102 131568 172170
rect 131248 172046 131318 172102
rect 131374 172046 131442 172102
rect 131498 172046 131568 172102
rect 131248 171978 131568 172046
rect 131248 171922 131318 171978
rect 131374 171922 131442 171978
rect 131498 171922 131568 171978
rect 131248 171888 131568 171922
rect 161968 172350 162288 172384
rect 161968 172294 162038 172350
rect 162094 172294 162162 172350
rect 162218 172294 162288 172350
rect 161968 172226 162288 172294
rect 161968 172170 162038 172226
rect 162094 172170 162162 172226
rect 162218 172170 162288 172226
rect 161968 172102 162288 172170
rect 161968 172046 162038 172102
rect 162094 172046 162162 172102
rect 162218 172046 162288 172102
rect 161968 171978 162288 172046
rect 161968 171922 162038 171978
rect 162094 171922 162162 171978
rect 162218 171922 162288 171978
rect 161968 171888 162288 171922
rect 192688 172350 193008 172384
rect 192688 172294 192758 172350
rect 192814 172294 192882 172350
rect 192938 172294 193008 172350
rect 192688 172226 193008 172294
rect 192688 172170 192758 172226
rect 192814 172170 192882 172226
rect 192938 172170 193008 172226
rect 192688 172102 193008 172170
rect 192688 172046 192758 172102
rect 192814 172046 192882 172102
rect 192938 172046 193008 172102
rect 192688 171978 193008 172046
rect 192688 171922 192758 171978
rect 192814 171922 192882 171978
rect 192938 171922 193008 171978
rect 192688 171888 193008 171922
rect 223408 172350 223728 172384
rect 223408 172294 223478 172350
rect 223534 172294 223602 172350
rect 223658 172294 223728 172350
rect 223408 172226 223728 172294
rect 223408 172170 223478 172226
rect 223534 172170 223602 172226
rect 223658 172170 223728 172226
rect 223408 172102 223728 172170
rect 223408 172046 223478 172102
rect 223534 172046 223602 172102
rect 223658 172046 223728 172102
rect 223408 171978 223728 172046
rect 223408 171922 223478 171978
rect 223534 171922 223602 171978
rect 223658 171922 223728 171978
rect 223408 171888 223728 171922
rect 254128 172350 254448 172384
rect 254128 172294 254198 172350
rect 254254 172294 254322 172350
rect 254378 172294 254448 172350
rect 254128 172226 254448 172294
rect 254128 172170 254198 172226
rect 254254 172170 254322 172226
rect 254378 172170 254448 172226
rect 254128 172102 254448 172170
rect 254128 172046 254198 172102
rect 254254 172046 254322 172102
rect 254378 172046 254448 172102
rect 254128 171978 254448 172046
rect 254128 171922 254198 171978
rect 254254 171922 254322 171978
rect 254378 171922 254448 171978
rect 254128 171888 254448 171922
rect 284848 172350 285168 172384
rect 284848 172294 284918 172350
rect 284974 172294 285042 172350
rect 285098 172294 285168 172350
rect 284848 172226 285168 172294
rect 284848 172170 284918 172226
rect 284974 172170 285042 172226
rect 285098 172170 285168 172226
rect 284848 172102 285168 172170
rect 284848 172046 284918 172102
rect 284974 172046 285042 172102
rect 285098 172046 285168 172102
rect 284848 171978 285168 172046
rect 284848 171922 284918 171978
rect 284974 171922 285042 171978
rect 285098 171922 285168 171978
rect 284848 171888 285168 171922
rect 315568 172350 315888 172384
rect 315568 172294 315638 172350
rect 315694 172294 315762 172350
rect 315818 172294 315888 172350
rect 315568 172226 315888 172294
rect 315568 172170 315638 172226
rect 315694 172170 315762 172226
rect 315818 172170 315888 172226
rect 315568 172102 315888 172170
rect 315568 172046 315638 172102
rect 315694 172046 315762 172102
rect 315818 172046 315888 172102
rect 315568 171978 315888 172046
rect 315568 171922 315638 171978
rect 315694 171922 315762 171978
rect 315818 171922 315888 171978
rect 315568 171888 315888 171922
rect 346288 172350 346608 172384
rect 346288 172294 346358 172350
rect 346414 172294 346482 172350
rect 346538 172294 346608 172350
rect 346288 172226 346608 172294
rect 346288 172170 346358 172226
rect 346414 172170 346482 172226
rect 346538 172170 346608 172226
rect 346288 172102 346608 172170
rect 346288 172046 346358 172102
rect 346414 172046 346482 172102
rect 346538 172046 346608 172102
rect 346288 171978 346608 172046
rect 346288 171922 346358 171978
rect 346414 171922 346482 171978
rect 346538 171922 346608 171978
rect 346288 171888 346608 171922
rect 377008 172350 377328 172384
rect 377008 172294 377078 172350
rect 377134 172294 377202 172350
rect 377258 172294 377328 172350
rect 377008 172226 377328 172294
rect 377008 172170 377078 172226
rect 377134 172170 377202 172226
rect 377258 172170 377328 172226
rect 377008 172102 377328 172170
rect 377008 172046 377078 172102
rect 377134 172046 377202 172102
rect 377258 172046 377328 172102
rect 377008 171978 377328 172046
rect 377008 171922 377078 171978
rect 377134 171922 377202 171978
rect 377258 171922 377328 171978
rect 377008 171888 377328 171922
rect 407728 172350 408048 172384
rect 407728 172294 407798 172350
rect 407854 172294 407922 172350
rect 407978 172294 408048 172350
rect 407728 172226 408048 172294
rect 407728 172170 407798 172226
rect 407854 172170 407922 172226
rect 407978 172170 408048 172226
rect 407728 172102 408048 172170
rect 407728 172046 407798 172102
rect 407854 172046 407922 172102
rect 407978 172046 408048 172102
rect 407728 171978 408048 172046
rect 407728 171922 407798 171978
rect 407854 171922 407922 171978
rect 407978 171922 408048 171978
rect 407728 171888 408048 171922
rect 438448 172350 438768 172384
rect 438448 172294 438518 172350
rect 438574 172294 438642 172350
rect 438698 172294 438768 172350
rect 438448 172226 438768 172294
rect 438448 172170 438518 172226
rect 438574 172170 438642 172226
rect 438698 172170 438768 172226
rect 438448 172102 438768 172170
rect 438448 172046 438518 172102
rect 438574 172046 438642 172102
rect 438698 172046 438768 172102
rect 438448 171978 438768 172046
rect 438448 171922 438518 171978
rect 438574 171922 438642 171978
rect 438698 171922 438768 171978
rect 438448 171888 438768 171922
rect 469168 172350 469488 172384
rect 469168 172294 469238 172350
rect 469294 172294 469362 172350
rect 469418 172294 469488 172350
rect 469168 172226 469488 172294
rect 469168 172170 469238 172226
rect 469294 172170 469362 172226
rect 469418 172170 469488 172226
rect 469168 172102 469488 172170
rect 469168 172046 469238 172102
rect 469294 172046 469362 172102
rect 469418 172046 469488 172102
rect 469168 171978 469488 172046
rect 469168 171922 469238 171978
rect 469294 171922 469362 171978
rect 469418 171922 469488 171978
rect 469168 171888 469488 171922
rect 499888 172350 500208 172384
rect 499888 172294 499958 172350
rect 500014 172294 500082 172350
rect 500138 172294 500208 172350
rect 499888 172226 500208 172294
rect 499888 172170 499958 172226
rect 500014 172170 500082 172226
rect 500138 172170 500208 172226
rect 499888 172102 500208 172170
rect 499888 172046 499958 172102
rect 500014 172046 500082 172102
rect 500138 172046 500208 172102
rect 499888 171978 500208 172046
rect 499888 171922 499958 171978
rect 500014 171922 500082 171978
rect 500138 171922 500208 171978
rect 499888 171888 500208 171922
rect 530608 172350 530928 172384
rect 530608 172294 530678 172350
rect 530734 172294 530802 172350
rect 530858 172294 530928 172350
rect 530608 172226 530928 172294
rect 530608 172170 530678 172226
rect 530734 172170 530802 172226
rect 530858 172170 530928 172226
rect 530608 172102 530928 172170
rect 530608 172046 530678 172102
rect 530734 172046 530802 172102
rect 530858 172046 530928 172102
rect 530608 171978 530928 172046
rect 530608 171922 530678 171978
rect 530734 171922 530802 171978
rect 530858 171922 530928 171978
rect 530608 171888 530928 171922
rect 111154 166294 111250 166350
rect 111306 166294 111374 166350
rect 111430 166294 111498 166350
rect 111554 166294 111622 166350
rect 111678 166294 111774 166350
rect 111154 166226 111774 166294
rect 111154 166170 111250 166226
rect 111306 166170 111374 166226
rect 111430 166170 111498 166226
rect 111554 166170 111622 166226
rect 111678 166170 111774 166226
rect 111154 166102 111774 166170
rect 111154 166046 111250 166102
rect 111306 166046 111374 166102
rect 111430 166046 111498 166102
rect 111554 166046 111622 166102
rect 111678 166046 111774 166102
rect 111154 165978 111774 166046
rect 111154 165922 111250 165978
rect 111306 165922 111374 165978
rect 111430 165922 111498 165978
rect 111554 165922 111622 165978
rect 111678 165922 111774 165978
rect 96874 154294 96970 154350
rect 97026 154294 97094 154350
rect 97150 154294 97218 154350
rect 97274 154294 97342 154350
rect 97398 154294 97494 154350
rect 96874 154226 97494 154294
rect 96874 154170 96970 154226
rect 97026 154170 97094 154226
rect 97150 154170 97218 154226
rect 97274 154170 97342 154226
rect 97398 154170 97494 154226
rect 96874 154102 97494 154170
rect 96874 154046 96970 154102
rect 97026 154046 97094 154102
rect 97150 154046 97218 154102
rect 97274 154046 97342 154102
rect 97398 154046 97494 154102
rect 96874 153978 97494 154046
rect 96874 153922 96970 153978
rect 97026 153922 97094 153978
rect 97150 153922 97218 153978
rect 97274 153922 97342 153978
rect 97398 153922 97494 153978
rect 96874 136350 97494 153922
rect 100528 154350 100848 154384
rect 100528 154294 100598 154350
rect 100654 154294 100722 154350
rect 100778 154294 100848 154350
rect 100528 154226 100848 154294
rect 100528 154170 100598 154226
rect 100654 154170 100722 154226
rect 100778 154170 100848 154226
rect 100528 154102 100848 154170
rect 100528 154046 100598 154102
rect 100654 154046 100722 154102
rect 100778 154046 100848 154102
rect 100528 153978 100848 154046
rect 100528 153922 100598 153978
rect 100654 153922 100722 153978
rect 100778 153922 100848 153978
rect 100528 153888 100848 153922
rect 111154 148350 111774 165922
rect 115888 166350 116208 166384
rect 115888 166294 115958 166350
rect 116014 166294 116082 166350
rect 116138 166294 116208 166350
rect 115888 166226 116208 166294
rect 115888 166170 115958 166226
rect 116014 166170 116082 166226
rect 116138 166170 116208 166226
rect 115888 166102 116208 166170
rect 115888 166046 115958 166102
rect 116014 166046 116082 166102
rect 116138 166046 116208 166102
rect 115888 165978 116208 166046
rect 115888 165922 115958 165978
rect 116014 165922 116082 165978
rect 116138 165922 116208 165978
rect 115888 165888 116208 165922
rect 146608 166350 146928 166384
rect 146608 166294 146678 166350
rect 146734 166294 146802 166350
rect 146858 166294 146928 166350
rect 146608 166226 146928 166294
rect 146608 166170 146678 166226
rect 146734 166170 146802 166226
rect 146858 166170 146928 166226
rect 146608 166102 146928 166170
rect 146608 166046 146678 166102
rect 146734 166046 146802 166102
rect 146858 166046 146928 166102
rect 146608 165978 146928 166046
rect 146608 165922 146678 165978
rect 146734 165922 146802 165978
rect 146858 165922 146928 165978
rect 146608 165888 146928 165922
rect 177328 166350 177648 166384
rect 177328 166294 177398 166350
rect 177454 166294 177522 166350
rect 177578 166294 177648 166350
rect 177328 166226 177648 166294
rect 177328 166170 177398 166226
rect 177454 166170 177522 166226
rect 177578 166170 177648 166226
rect 177328 166102 177648 166170
rect 177328 166046 177398 166102
rect 177454 166046 177522 166102
rect 177578 166046 177648 166102
rect 177328 165978 177648 166046
rect 177328 165922 177398 165978
rect 177454 165922 177522 165978
rect 177578 165922 177648 165978
rect 177328 165888 177648 165922
rect 208048 166350 208368 166384
rect 208048 166294 208118 166350
rect 208174 166294 208242 166350
rect 208298 166294 208368 166350
rect 208048 166226 208368 166294
rect 208048 166170 208118 166226
rect 208174 166170 208242 166226
rect 208298 166170 208368 166226
rect 208048 166102 208368 166170
rect 208048 166046 208118 166102
rect 208174 166046 208242 166102
rect 208298 166046 208368 166102
rect 208048 165978 208368 166046
rect 208048 165922 208118 165978
rect 208174 165922 208242 165978
rect 208298 165922 208368 165978
rect 208048 165888 208368 165922
rect 238768 166350 239088 166384
rect 238768 166294 238838 166350
rect 238894 166294 238962 166350
rect 239018 166294 239088 166350
rect 238768 166226 239088 166294
rect 238768 166170 238838 166226
rect 238894 166170 238962 166226
rect 239018 166170 239088 166226
rect 238768 166102 239088 166170
rect 238768 166046 238838 166102
rect 238894 166046 238962 166102
rect 239018 166046 239088 166102
rect 238768 165978 239088 166046
rect 238768 165922 238838 165978
rect 238894 165922 238962 165978
rect 239018 165922 239088 165978
rect 238768 165888 239088 165922
rect 269488 166350 269808 166384
rect 269488 166294 269558 166350
rect 269614 166294 269682 166350
rect 269738 166294 269808 166350
rect 269488 166226 269808 166294
rect 269488 166170 269558 166226
rect 269614 166170 269682 166226
rect 269738 166170 269808 166226
rect 269488 166102 269808 166170
rect 269488 166046 269558 166102
rect 269614 166046 269682 166102
rect 269738 166046 269808 166102
rect 269488 165978 269808 166046
rect 269488 165922 269558 165978
rect 269614 165922 269682 165978
rect 269738 165922 269808 165978
rect 269488 165888 269808 165922
rect 300208 166350 300528 166384
rect 300208 166294 300278 166350
rect 300334 166294 300402 166350
rect 300458 166294 300528 166350
rect 300208 166226 300528 166294
rect 300208 166170 300278 166226
rect 300334 166170 300402 166226
rect 300458 166170 300528 166226
rect 300208 166102 300528 166170
rect 300208 166046 300278 166102
rect 300334 166046 300402 166102
rect 300458 166046 300528 166102
rect 300208 165978 300528 166046
rect 300208 165922 300278 165978
rect 300334 165922 300402 165978
rect 300458 165922 300528 165978
rect 300208 165888 300528 165922
rect 330928 166350 331248 166384
rect 330928 166294 330998 166350
rect 331054 166294 331122 166350
rect 331178 166294 331248 166350
rect 330928 166226 331248 166294
rect 330928 166170 330998 166226
rect 331054 166170 331122 166226
rect 331178 166170 331248 166226
rect 330928 166102 331248 166170
rect 330928 166046 330998 166102
rect 331054 166046 331122 166102
rect 331178 166046 331248 166102
rect 330928 165978 331248 166046
rect 330928 165922 330998 165978
rect 331054 165922 331122 165978
rect 331178 165922 331248 165978
rect 330928 165888 331248 165922
rect 361648 166350 361968 166384
rect 361648 166294 361718 166350
rect 361774 166294 361842 166350
rect 361898 166294 361968 166350
rect 361648 166226 361968 166294
rect 361648 166170 361718 166226
rect 361774 166170 361842 166226
rect 361898 166170 361968 166226
rect 361648 166102 361968 166170
rect 361648 166046 361718 166102
rect 361774 166046 361842 166102
rect 361898 166046 361968 166102
rect 361648 165978 361968 166046
rect 361648 165922 361718 165978
rect 361774 165922 361842 165978
rect 361898 165922 361968 165978
rect 361648 165888 361968 165922
rect 392368 166350 392688 166384
rect 392368 166294 392438 166350
rect 392494 166294 392562 166350
rect 392618 166294 392688 166350
rect 392368 166226 392688 166294
rect 392368 166170 392438 166226
rect 392494 166170 392562 166226
rect 392618 166170 392688 166226
rect 392368 166102 392688 166170
rect 392368 166046 392438 166102
rect 392494 166046 392562 166102
rect 392618 166046 392688 166102
rect 392368 165978 392688 166046
rect 392368 165922 392438 165978
rect 392494 165922 392562 165978
rect 392618 165922 392688 165978
rect 392368 165888 392688 165922
rect 423088 166350 423408 166384
rect 423088 166294 423158 166350
rect 423214 166294 423282 166350
rect 423338 166294 423408 166350
rect 423088 166226 423408 166294
rect 423088 166170 423158 166226
rect 423214 166170 423282 166226
rect 423338 166170 423408 166226
rect 423088 166102 423408 166170
rect 423088 166046 423158 166102
rect 423214 166046 423282 166102
rect 423338 166046 423408 166102
rect 423088 165978 423408 166046
rect 423088 165922 423158 165978
rect 423214 165922 423282 165978
rect 423338 165922 423408 165978
rect 423088 165888 423408 165922
rect 453808 166350 454128 166384
rect 453808 166294 453878 166350
rect 453934 166294 454002 166350
rect 454058 166294 454128 166350
rect 453808 166226 454128 166294
rect 453808 166170 453878 166226
rect 453934 166170 454002 166226
rect 454058 166170 454128 166226
rect 453808 166102 454128 166170
rect 453808 166046 453878 166102
rect 453934 166046 454002 166102
rect 454058 166046 454128 166102
rect 453808 165978 454128 166046
rect 453808 165922 453878 165978
rect 453934 165922 454002 165978
rect 454058 165922 454128 165978
rect 453808 165888 454128 165922
rect 484528 166350 484848 166384
rect 484528 166294 484598 166350
rect 484654 166294 484722 166350
rect 484778 166294 484848 166350
rect 484528 166226 484848 166294
rect 484528 166170 484598 166226
rect 484654 166170 484722 166226
rect 484778 166170 484848 166226
rect 484528 166102 484848 166170
rect 484528 166046 484598 166102
rect 484654 166046 484722 166102
rect 484778 166046 484848 166102
rect 484528 165978 484848 166046
rect 484528 165922 484598 165978
rect 484654 165922 484722 165978
rect 484778 165922 484848 165978
rect 484528 165888 484848 165922
rect 515248 166350 515568 166384
rect 515248 166294 515318 166350
rect 515374 166294 515442 166350
rect 515498 166294 515568 166350
rect 515248 166226 515568 166294
rect 515248 166170 515318 166226
rect 515374 166170 515442 166226
rect 515498 166170 515568 166226
rect 515248 166102 515568 166170
rect 515248 166046 515318 166102
rect 515374 166046 515442 166102
rect 515498 166046 515568 166102
rect 515248 165978 515568 166046
rect 515248 165922 515318 165978
rect 515374 165922 515442 165978
rect 515498 165922 515568 165978
rect 515248 165888 515568 165922
rect 545968 166350 546288 166384
rect 545968 166294 546038 166350
rect 546094 166294 546162 166350
rect 546218 166294 546288 166350
rect 545968 166226 546288 166294
rect 545968 166170 546038 166226
rect 546094 166170 546162 166226
rect 546218 166170 546288 166226
rect 545968 166102 546288 166170
rect 545968 166046 546038 166102
rect 546094 166046 546162 166102
rect 546218 166046 546288 166102
rect 545968 165978 546288 166046
rect 545968 165922 546038 165978
rect 546094 165922 546162 165978
rect 546218 165922 546288 165978
rect 545968 165888 546288 165922
rect 561154 166350 561774 183922
rect 561154 166294 561250 166350
rect 561306 166294 561374 166350
rect 561430 166294 561498 166350
rect 561554 166294 561622 166350
rect 561678 166294 561774 166350
rect 561154 166226 561774 166294
rect 561154 166170 561250 166226
rect 561306 166170 561374 166226
rect 561430 166170 561498 166226
rect 561554 166170 561622 166226
rect 561678 166170 561774 166226
rect 561154 166102 561774 166170
rect 561154 166046 561250 166102
rect 561306 166046 561374 166102
rect 561430 166046 561498 166102
rect 561554 166046 561622 166102
rect 561678 166046 561774 166102
rect 561154 165978 561774 166046
rect 561154 165922 561250 165978
rect 561306 165922 561374 165978
rect 561430 165922 561498 165978
rect 561554 165922 561622 165978
rect 561678 165922 561774 165978
rect 131248 154350 131568 154384
rect 131248 154294 131318 154350
rect 131374 154294 131442 154350
rect 131498 154294 131568 154350
rect 131248 154226 131568 154294
rect 131248 154170 131318 154226
rect 131374 154170 131442 154226
rect 131498 154170 131568 154226
rect 131248 154102 131568 154170
rect 131248 154046 131318 154102
rect 131374 154046 131442 154102
rect 131498 154046 131568 154102
rect 131248 153978 131568 154046
rect 131248 153922 131318 153978
rect 131374 153922 131442 153978
rect 131498 153922 131568 153978
rect 131248 153888 131568 153922
rect 161968 154350 162288 154384
rect 161968 154294 162038 154350
rect 162094 154294 162162 154350
rect 162218 154294 162288 154350
rect 161968 154226 162288 154294
rect 161968 154170 162038 154226
rect 162094 154170 162162 154226
rect 162218 154170 162288 154226
rect 161968 154102 162288 154170
rect 161968 154046 162038 154102
rect 162094 154046 162162 154102
rect 162218 154046 162288 154102
rect 161968 153978 162288 154046
rect 161968 153922 162038 153978
rect 162094 153922 162162 153978
rect 162218 153922 162288 153978
rect 161968 153888 162288 153922
rect 192688 154350 193008 154384
rect 192688 154294 192758 154350
rect 192814 154294 192882 154350
rect 192938 154294 193008 154350
rect 192688 154226 193008 154294
rect 192688 154170 192758 154226
rect 192814 154170 192882 154226
rect 192938 154170 193008 154226
rect 192688 154102 193008 154170
rect 192688 154046 192758 154102
rect 192814 154046 192882 154102
rect 192938 154046 193008 154102
rect 192688 153978 193008 154046
rect 192688 153922 192758 153978
rect 192814 153922 192882 153978
rect 192938 153922 193008 153978
rect 192688 153888 193008 153922
rect 223408 154350 223728 154384
rect 223408 154294 223478 154350
rect 223534 154294 223602 154350
rect 223658 154294 223728 154350
rect 223408 154226 223728 154294
rect 223408 154170 223478 154226
rect 223534 154170 223602 154226
rect 223658 154170 223728 154226
rect 223408 154102 223728 154170
rect 223408 154046 223478 154102
rect 223534 154046 223602 154102
rect 223658 154046 223728 154102
rect 223408 153978 223728 154046
rect 223408 153922 223478 153978
rect 223534 153922 223602 153978
rect 223658 153922 223728 153978
rect 223408 153888 223728 153922
rect 254128 154350 254448 154384
rect 254128 154294 254198 154350
rect 254254 154294 254322 154350
rect 254378 154294 254448 154350
rect 254128 154226 254448 154294
rect 254128 154170 254198 154226
rect 254254 154170 254322 154226
rect 254378 154170 254448 154226
rect 254128 154102 254448 154170
rect 254128 154046 254198 154102
rect 254254 154046 254322 154102
rect 254378 154046 254448 154102
rect 254128 153978 254448 154046
rect 254128 153922 254198 153978
rect 254254 153922 254322 153978
rect 254378 153922 254448 153978
rect 254128 153888 254448 153922
rect 284848 154350 285168 154384
rect 284848 154294 284918 154350
rect 284974 154294 285042 154350
rect 285098 154294 285168 154350
rect 284848 154226 285168 154294
rect 284848 154170 284918 154226
rect 284974 154170 285042 154226
rect 285098 154170 285168 154226
rect 284848 154102 285168 154170
rect 284848 154046 284918 154102
rect 284974 154046 285042 154102
rect 285098 154046 285168 154102
rect 284848 153978 285168 154046
rect 284848 153922 284918 153978
rect 284974 153922 285042 153978
rect 285098 153922 285168 153978
rect 284848 153888 285168 153922
rect 315568 154350 315888 154384
rect 315568 154294 315638 154350
rect 315694 154294 315762 154350
rect 315818 154294 315888 154350
rect 315568 154226 315888 154294
rect 315568 154170 315638 154226
rect 315694 154170 315762 154226
rect 315818 154170 315888 154226
rect 315568 154102 315888 154170
rect 315568 154046 315638 154102
rect 315694 154046 315762 154102
rect 315818 154046 315888 154102
rect 315568 153978 315888 154046
rect 315568 153922 315638 153978
rect 315694 153922 315762 153978
rect 315818 153922 315888 153978
rect 315568 153888 315888 153922
rect 346288 154350 346608 154384
rect 346288 154294 346358 154350
rect 346414 154294 346482 154350
rect 346538 154294 346608 154350
rect 346288 154226 346608 154294
rect 346288 154170 346358 154226
rect 346414 154170 346482 154226
rect 346538 154170 346608 154226
rect 346288 154102 346608 154170
rect 346288 154046 346358 154102
rect 346414 154046 346482 154102
rect 346538 154046 346608 154102
rect 346288 153978 346608 154046
rect 346288 153922 346358 153978
rect 346414 153922 346482 153978
rect 346538 153922 346608 153978
rect 346288 153888 346608 153922
rect 377008 154350 377328 154384
rect 377008 154294 377078 154350
rect 377134 154294 377202 154350
rect 377258 154294 377328 154350
rect 377008 154226 377328 154294
rect 377008 154170 377078 154226
rect 377134 154170 377202 154226
rect 377258 154170 377328 154226
rect 377008 154102 377328 154170
rect 377008 154046 377078 154102
rect 377134 154046 377202 154102
rect 377258 154046 377328 154102
rect 377008 153978 377328 154046
rect 377008 153922 377078 153978
rect 377134 153922 377202 153978
rect 377258 153922 377328 153978
rect 377008 153888 377328 153922
rect 407728 154350 408048 154384
rect 407728 154294 407798 154350
rect 407854 154294 407922 154350
rect 407978 154294 408048 154350
rect 407728 154226 408048 154294
rect 407728 154170 407798 154226
rect 407854 154170 407922 154226
rect 407978 154170 408048 154226
rect 407728 154102 408048 154170
rect 407728 154046 407798 154102
rect 407854 154046 407922 154102
rect 407978 154046 408048 154102
rect 407728 153978 408048 154046
rect 407728 153922 407798 153978
rect 407854 153922 407922 153978
rect 407978 153922 408048 153978
rect 407728 153888 408048 153922
rect 438448 154350 438768 154384
rect 438448 154294 438518 154350
rect 438574 154294 438642 154350
rect 438698 154294 438768 154350
rect 438448 154226 438768 154294
rect 438448 154170 438518 154226
rect 438574 154170 438642 154226
rect 438698 154170 438768 154226
rect 438448 154102 438768 154170
rect 438448 154046 438518 154102
rect 438574 154046 438642 154102
rect 438698 154046 438768 154102
rect 438448 153978 438768 154046
rect 438448 153922 438518 153978
rect 438574 153922 438642 153978
rect 438698 153922 438768 153978
rect 438448 153888 438768 153922
rect 469168 154350 469488 154384
rect 469168 154294 469238 154350
rect 469294 154294 469362 154350
rect 469418 154294 469488 154350
rect 469168 154226 469488 154294
rect 469168 154170 469238 154226
rect 469294 154170 469362 154226
rect 469418 154170 469488 154226
rect 469168 154102 469488 154170
rect 469168 154046 469238 154102
rect 469294 154046 469362 154102
rect 469418 154046 469488 154102
rect 469168 153978 469488 154046
rect 469168 153922 469238 153978
rect 469294 153922 469362 153978
rect 469418 153922 469488 153978
rect 469168 153888 469488 153922
rect 499888 154350 500208 154384
rect 499888 154294 499958 154350
rect 500014 154294 500082 154350
rect 500138 154294 500208 154350
rect 499888 154226 500208 154294
rect 499888 154170 499958 154226
rect 500014 154170 500082 154226
rect 500138 154170 500208 154226
rect 499888 154102 500208 154170
rect 499888 154046 499958 154102
rect 500014 154046 500082 154102
rect 500138 154046 500208 154102
rect 499888 153978 500208 154046
rect 499888 153922 499958 153978
rect 500014 153922 500082 153978
rect 500138 153922 500208 153978
rect 499888 153888 500208 153922
rect 530608 154350 530928 154384
rect 530608 154294 530678 154350
rect 530734 154294 530802 154350
rect 530858 154294 530928 154350
rect 530608 154226 530928 154294
rect 530608 154170 530678 154226
rect 530734 154170 530802 154226
rect 530858 154170 530928 154226
rect 530608 154102 530928 154170
rect 530608 154046 530678 154102
rect 530734 154046 530802 154102
rect 530858 154046 530928 154102
rect 530608 153978 530928 154046
rect 530608 153922 530678 153978
rect 530734 153922 530802 153978
rect 530858 153922 530928 153978
rect 530608 153888 530928 153922
rect 111154 148294 111250 148350
rect 111306 148294 111374 148350
rect 111430 148294 111498 148350
rect 111554 148294 111622 148350
rect 111678 148294 111774 148350
rect 111154 148226 111774 148294
rect 111154 148170 111250 148226
rect 111306 148170 111374 148226
rect 111430 148170 111498 148226
rect 111554 148170 111622 148226
rect 111678 148170 111774 148226
rect 111154 148102 111774 148170
rect 111154 148046 111250 148102
rect 111306 148046 111374 148102
rect 111430 148046 111498 148102
rect 111554 148046 111622 148102
rect 111678 148046 111774 148102
rect 111154 147978 111774 148046
rect 111154 147922 111250 147978
rect 111306 147922 111374 147978
rect 111430 147922 111498 147978
rect 111554 147922 111622 147978
rect 111678 147922 111774 147978
rect 96874 136294 96970 136350
rect 97026 136294 97094 136350
rect 97150 136294 97218 136350
rect 97274 136294 97342 136350
rect 97398 136294 97494 136350
rect 96874 136226 97494 136294
rect 96874 136170 96970 136226
rect 97026 136170 97094 136226
rect 97150 136170 97218 136226
rect 97274 136170 97342 136226
rect 97398 136170 97494 136226
rect 96874 136102 97494 136170
rect 96874 136046 96970 136102
rect 97026 136046 97094 136102
rect 97150 136046 97218 136102
rect 97274 136046 97342 136102
rect 97398 136046 97494 136102
rect 96874 135978 97494 136046
rect 96874 135922 96970 135978
rect 97026 135922 97094 135978
rect 97150 135922 97218 135978
rect 97274 135922 97342 135978
rect 97398 135922 97494 135978
rect 96874 118350 97494 135922
rect 100528 136350 100848 136384
rect 100528 136294 100598 136350
rect 100654 136294 100722 136350
rect 100778 136294 100848 136350
rect 100528 136226 100848 136294
rect 100528 136170 100598 136226
rect 100654 136170 100722 136226
rect 100778 136170 100848 136226
rect 100528 136102 100848 136170
rect 100528 136046 100598 136102
rect 100654 136046 100722 136102
rect 100778 136046 100848 136102
rect 100528 135978 100848 136046
rect 100528 135922 100598 135978
rect 100654 135922 100722 135978
rect 100778 135922 100848 135978
rect 100528 135888 100848 135922
rect 111154 130350 111774 147922
rect 115888 148350 116208 148384
rect 115888 148294 115958 148350
rect 116014 148294 116082 148350
rect 116138 148294 116208 148350
rect 115888 148226 116208 148294
rect 115888 148170 115958 148226
rect 116014 148170 116082 148226
rect 116138 148170 116208 148226
rect 115888 148102 116208 148170
rect 115888 148046 115958 148102
rect 116014 148046 116082 148102
rect 116138 148046 116208 148102
rect 115888 147978 116208 148046
rect 115888 147922 115958 147978
rect 116014 147922 116082 147978
rect 116138 147922 116208 147978
rect 115888 147888 116208 147922
rect 146608 148350 146928 148384
rect 146608 148294 146678 148350
rect 146734 148294 146802 148350
rect 146858 148294 146928 148350
rect 146608 148226 146928 148294
rect 146608 148170 146678 148226
rect 146734 148170 146802 148226
rect 146858 148170 146928 148226
rect 146608 148102 146928 148170
rect 146608 148046 146678 148102
rect 146734 148046 146802 148102
rect 146858 148046 146928 148102
rect 146608 147978 146928 148046
rect 146608 147922 146678 147978
rect 146734 147922 146802 147978
rect 146858 147922 146928 147978
rect 146608 147888 146928 147922
rect 177328 148350 177648 148384
rect 177328 148294 177398 148350
rect 177454 148294 177522 148350
rect 177578 148294 177648 148350
rect 177328 148226 177648 148294
rect 177328 148170 177398 148226
rect 177454 148170 177522 148226
rect 177578 148170 177648 148226
rect 177328 148102 177648 148170
rect 177328 148046 177398 148102
rect 177454 148046 177522 148102
rect 177578 148046 177648 148102
rect 177328 147978 177648 148046
rect 177328 147922 177398 147978
rect 177454 147922 177522 147978
rect 177578 147922 177648 147978
rect 177328 147888 177648 147922
rect 208048 148350 208368 148384
rect 208048 148294 208118 148350
rect 208174 148294 208242 148350
rect 208298 148294 208368 148350
rect 208048 148226 208368 148294
rect 208048 148170 208118 148226
rect 208174 148170 208242 148226
rect 208298 148170 208368 148226
rect 208048 148102 208368 148170
rect 208048 148046 208118 148102
rect 208174 148046 208242 148102
rect 208298 148046 208368 148102
rect 208048 147978 208368 148046
rect 208048 147922 208118 147978
rect 208174 147922 208242 147978
rect 208298 147922 208368 147978
rect 208048 147888 208368 147922
rect 238768 148350 239088 148384
rect 238768 148294 238838 148350
rect 238894 148294 238962 148350
rect 239018 148294 239088 148350
rect 238768 148226 239088 148294
rect 238768 148170 238838 148226
rect 238894 148170 238962 148226
rect 239018 148170 239088 148226
rect 238768 148102 239088 148170
rect 238768 148046 238838 148102
rect 238894 148046 238962 148102
rect 239018 148046 239088 148102
rect 238768 147978 239088 148046
rect 238768 147922 238838 147978
rect 238894 147922 238962 147978
rect 239018 147922 239088 147978
rect 238768 147888 239088 147922
rect 269488 148350 269808 148384
rect 269488 148294 269558 148350
rect 269614 148294 269682 148350
rect 269738 148294 269808 148350
rect 269488 148226 269808 148294
rect 269488 148170 269558 148226
rect 269614 148170 269682 148226
rect 269738 148170 269808 148226
rect 269488 148102 269808 148170
rect 269488 148046 269558 148102
rect 269614 148046 269682 148102
rect 269738 148046 269808 148102
rect 269488 147978 269808 148046
rect 269488 147922 269558 147978
rect 269614 147922 269682 147978
rect 269738 147922 269808 147978
rect 269488 147888 269808 147922
rect 300208 148350 300528 148384
rect 300208 148294 300278 148350
rect 300334 148294 300402 148350
rect 300458 148294 300528 148350
rect 300208 148226 300528 148294
rect 300208 148170 300278 148226
rect 300334 148170 300402 148226
rect 300458 148170 300528 148226
rect 300208 148102 300528 148170
rect 300208 148046 300278 148102
rect 300334 148046 300402 148102
rect 300458 148046 300528 148102
rect 300208 147978 300528 148046
rect 300208 147922 300278 147978
rect 300334 147922 300402 147978
rect 300458 147922 300528 147978
rect 300208 147888 300528 147922
rect 330928 148350 331248 148384
rect 330928 148294 330998 148350
rect 331054 148294 331122 148350
rect 331178 148294 331248 148350
rect 330928 148226 331248 148294
rect 330928 148170 330998 148226
rect 331054 148170 331122 148226
rect 331178 148170 331248 148226
rect 330928 148102 331248 148170
rect 330928 148046 330998 148102
rect 331054 148046 331122 148102
rect 331178 148046 331248 148102
rect 330928 147978 331248 148046
rect 330928 147922 330998 147978
rect 331054 147922 331122 147978
rect 331178 147922 331248 147978
rect 330928 147888 331248 147922
rect 361648 148350 361968 148384
rect 361648 148294 361718 148350
rect 361774 148294 361842 148350
rect 361898 148294 361968 148350
rect 361648 148226 361968 148294
rect 361648 148170 361718 148226
rect 361774 148170 361842 148226
rect 361898 148170 361968 148226
rect 361648 148102 361968 148170
rect 361648 148046 361718 148102
rect 361774 148046 361842 148102
rect 361898 148046 361968 148102
rect 361648 147978 361968 148046
rect 361648 147922 361718 147978
rect 361774 147922 361842 147978
rect 361898 147922 361968 147978
rect 361648 147888 361968 147922
rect 392368 148350 392688 148384
rect 392368 148294 392438 148350
rect 392494 148294 392562 148350
rect 392618 148294 392688 148350
rect 392368 148226 392688 148294
rect 392368 148170 392438 148226
rect 392494 148170 392562 148226
rect 392618 148170 392688 148226
rect 392368 148102 392688 148170
rect 392368 148046 392438 148102
rect 392494 148046 392562 148102
rect 392618 148046 392688 148102
rect 392368 147978 392688 148046
rect 392368 147922 392438 147978
rect 392494 147922 392562 147978
rect 392618 147922 392688 147978
rect 392368 147888 392688 147922
rect 423088 148350 423408 148384
rect 423088 148294 423158 148350
rect 423214 148294 423282 148350
rect 423338 148294 423408 148350
rect 423088 148226 423408 148294
rect 423088 148170 423158 148226
rect 423214 148170 423282 148226
rect 423338 148170 423408 148226
rect 423088 148102 423408 148170
rect 423088 148046 423158 148102
rect 423214 148046 423282 148102
rect 423338 148046 423408 148102
rect 423088 147978 423408 148046
rect 423088 147922 423158 147978
rect 423214 147922 423282 147978
rect 423338 147922 423408 147978
rect 423088 147888 423408 147922
rect 453808 148350 454128 148384
rect 453808 148294 453878 148350
rect 453934 148294 454002 148350
rect 454058 148294 454128 148350
rect 453808 148226 454128 148294
rect 453808 148170 453878 148226
rect 453934 148170 454002 148226
rect 454058 148170 454128 148226
rect 453808 148102 454128 148170
rect 453808 148046 453878 148102
rect 453934 148046 454002 148102
rect 454058 148046 454128 148102
rect 453808 147978 454128 148046
rect 453808 147922 453878 147978
rect 453934 147922 454002 147978
rect 454058 147922 454128 147978
rect 453808 147888 454128 147922
rect 484528 148350 484848 148384
rect 484528 148294 484598 148350
rect 484654 148294 484722 148350
rect 484778 148294 484848 148350
rect 484528 148226 484848 148294
rect 484528 148170 484598 148226
rect 484654 148170 484722 148226
rect 484778 148170 484848 148226
rect 484528 148102 484848 148170
rect 484528 148046 484598 148102
rect 484654 148046 484722 148102
rect 484778 148046 484848 148102
rect 484528 147978 484848 148046
rect 484528 147922 484598 147978
rect 484654 147922 484722 147978
rect 484778 147922 484848 147978
rect 484528 147888 484848 147922
rect 515248 148350 515568 148384
rect 515248 148294 515318 148350
rect 515374 148294 515442 148350
rect 515498 148294 515568 148350
rect 515248 148226 515568 148294
rect 515248 148170 515318 148226
rect 515374 148170 515442 148226
rect 515498 148170 515568 148226
rect 515248 148102 515568 148170
rect 515248 148046 515318 148102
rect 515374 148046 515442 148102
rect 515498 148046 515568 148102
rect 515248 147978 515568 148046
rect 515248 147922 515318 147978
rect 515374 147922 515442 147978
rect 515498 147922 515568 147978
rect 515248 147888 515568 147922
rect 545968 148350 546288 148384
rect 545968 148294 546038 148350
rect 546094 148294 546162 148350
rect 546218 148294 546288 148350
rect 545968 148226 546288 148294
rect 545968 148170 546038 148226
rect 546094 148170 546162 148226
rect 546218 148170 546288 148226
rect 545968 148102 546288 148170
rect 545968 148046 546038 148102
rect 546094 148046 546162 148102
rect 546218 148046 546288 148102
rect 545968 147978 546288 148046
rect 545968 147922 546038 147978
rect 546094 147922 546162 147978
rect 546218 147922 546288 147978
rect 545968 147888 546288 147922
rect 561154 148350 561774 165922
rect 561154 148294 561250 148350
rect 561306 148294 561374 148350
rect 561430 148294 561498 148350
rect 561554 148294 561622 148350
rect 561678 148294 561774 148350
rect 561154 148226 561774 148294
rect 561154 148170 561250 148226
rect 561306 148170 561374 148226
rect 561430 148170 561498 148226
rect 561554 148170 561622 148226
rect 561678 148170 561774 148226
rect 561154 148102 561774 148170
rect 561154 148046 561250 148102
rect 561306 148046 561374 148102
rect 561430 148046 561498 148102
rect 561554 148046 561622 148102
rect 561678 148046 561774 148102
rect 561154 147978 561774 148046
rect 561154 147922 561250 147978
rect 561306 147922 561374 147978
rect 561430 147922 561498 147978
rect 561554 147922 561622 147978
rect 561678 147922 561774 147978
rect 131248 136350 131568 136384
rect 131248 136294 131318 136350
rect 131374 136294 131442 136350
rect 131498 136294 131568 136350
rect 131248 136226 131568 136294
rect 131248 136170 131318 136226
rect 131374 136170 131442 136226
rect 131498 136170 131568 136226
rect 131248 136102 131568 136170
rect 131248 136046 131318 136102
rect 131374 136046 131442 136102
rect 131498 136046 131568 136102
rect 131248 135978 131568 136046
rect 131248 135922 131318 135978
rect 131374 135922 131442 135978
rect 131498 135922 131568 135978
rect 131248 135888 131568 135922
rect 161968 136350 162288 136384
rect 161968 136294 162038 136350
rect 162094 136294 162162 136350
rect 162218 136294 162288 136350
rect 161968 136226 162288 136294
rect 161968 136170 162038 136226
rect 162094 136170 162162 136226
rect 162218 136170 162288 136226
rect 161968 136102 162288 136170
rect 161968 136046 162038 136102
rect 162094 136046 162162 136102
rect 162218 136046 162288 136102
rect 161968 135978 162288 136046
rect 161968 135922 162038 135978
rect 162094 135922 162162 135978
rect 162218 135922 162288 135978
rect 161968 135888 162288 135922
rect 192688 136350 193008 136384
rect 192688 136294 192758 136350
rect 192814 136294 192882 136350
rect 192938 136294 193008 136350
rect 192688 136226 193008 136294
rect 192688 136170 192758 136226
rect 192814 136170 192882 136226
rect 192938 136170 193008 136226
rect 192688 136102 193008 136170
rect 192688 136046 192758 136102
rect 192814 136046 192882 136102
rect 192938 136046 193008 136102
rect 192688 135978 193008 136046
rect 192688 135922 192758 135978
rect 192814 135922 192882 135978
rect 192938 135922 193008 135978
rect 192688 135888 193008 135922
rect 223408 136350 223728 136384
rect 223408 136294 223478 136350
rect 223534 136294 223602 136350
rect 223658 136294 223728 136350
rect 223408 136226 223728 136294
rect 223408 136170 223478 136226
rect 223534 136170 223602 136226
rect 223658 136170 223728 136226
rect 223408 136102 223728 136170
rect 223408 136046 223478 136102
rect 223534 136046 223602 136102
rect 223658 136046 223728 136102
rect 223408 135978 223728 136046
rect 223408 135922 223478 135978
rect 223534 135922 223602 135978
rect 223658 135922 223728 135978
rect 223408 135888 223728 135922
rect 254128 136350 254448 136384
rect 254128 136294 254198 136350
rect 254254 136294 254322 136350
rect 254378 136294 254448 136350
rect 254128 136226 254448 136294
rect 254128 136170 254198 136226
rect 254254 136170 254322 136226
rect 254378 136170 254448 136226
rect 254128 136102 254448 136170
rect 254128 136046 254198 136102
rect 254254 136046 254322 136102
rect 254378 136046 254448 136102
rect 254128 135978 254448 136046
rect 254128 135922 254198 135978
rect 254254 135922 254322 135978
rect 254378 135922 254448 135978
rect 254128 135888 254448 135922
rect 284848 136350 285168 136384
rect 284848 136294 284918 136350
rect 284974 136294 285042 136350
rect 285098 136294 285168 136350
rect 284848 136226 285168 136294
rect 284848 136170 284918 136226
rect 284974 136170 285042 136226
rect 285098 136170 285168 136226
rect 284848 136102 285168 136170
rect 284848 136046 284918 136102
rect 284974 136046 285042 136102
rect 285098 136046 285168 136102
rect 284848 135978 285168 136046
rect 284848 135922 284918 135978
rect 284974 135922 285042 135978
rect 285098 135922 285168 135978
rect 284848 135888 285168 135922
rect 315568 136350 315888 136384
rect 315568 136294 315638 136350
rect 315694 136294 315762 136350
rect 315818 136294 315888 136350
rect 315568 136226 315888 136294
rect 315568 136170 315638 136226
rect 315694 136170 315762 136226
rect 315818 136170 315888 136226
rect 315568 136102 315888 136170
rect 315568 136046 315638 136102
rect 315694 136046 315762 136102
rect 315818 136046 315888 136102
rect 315568 135978 315888 136046
rect 315568 135922 315638 135978
rect 315694 135922 315762 135978
rect 315818 135922 315888 135978
rect 315568 135888 315888 135922
rect 346288 136350 346608 136384
rect 346288 136294 346358 136350
rect 346414 136294 346482 136350
rect 346538 136294 346608 136350
rect 346288 136226 346608 136294
rect 346288 136170 346358 136226
rect 346414 136170 346482 136226
rect 346538 136170 346608 136226
rect 346288 136102 346608 136170
rect 346288 136046 346358 136102
rect 346414 136046 346482 136102
rect 346538 136046 346608 136102
rect 346288 135978 346608 136046
rect 346288 135922 346358 135978
rect 346414 135922 346482 135978
rect 346538 135922 346608 135978
rect 346288 135888 346608 135922
rect 377008 136350 377328 136384
rect 377008 136294 377078 136350
rect 377134 136294 377202 136350
rect 377258 136294 377328 136350
rect 377008 136226 377328 136294
rect 377008 136170 377078 136226
rect 377134 136170 377202 136226
rect 377258 136170 377328 136226
rect 377008 136102 377328 136170
rect 377008 136046 377078 136102
rect 377134 136046 377202 136102
rect 377258 136046 377328 136102
rect 377008 135978 377328 136046
rect 377008 135922 377078 135978
rect 377134 135922 377202 135978
rect 377258 135922 377328 135978
rect 377008 135888 377328 135922
rect 407728 136350 408048 136384
rect 407728 136294 407798 136350
rect 407854 136294 407922 136350
rect 407978 136294 408048 136350
rect 407728 136226 408048 136294
rect 407728 136170 407798 136226
rect 407854 136170 407922 136226
rect 407978 136170 408048 136226
rect 407728 136102 408048 136170
rect 407728 136046 407798 136102
rect 407854 136046 407922 136102
rect 407978 136046 408048 136102
rect 407728 135978 408048 136046
rect 407728 135922 407798 135978
rect 407854 135922 407922 135978
rect 407978 135922 408048 135978
rect 407728 135888 408048 135922
rect 438448 136350 438768 136384
rect 438448 136294 438518 136350
rect 438574 136294 438642 136350
rect 438698 136294 438768 136350
rect 438448 136226 438768 136294
rect 438448 136170 438518 136226
rect 438574 136170 438642 136226
rect 438698 136170 438768 136226
rect 438448 136102 438768 136170
rect 438448 136046 438518 136102
rect 438574 136046 438642 136102
rect 438698 136046 438768 136102
rect 438448 135978 438768 136046
rect 438448 135922 438518 135978
rect 438574 135922 438642 135978
rect 438698 135922 438768 135978
rect 438448 135888 438768 135922
rect 469168 136350 469488 136384
rect 469168 136294 469238 136350
rect 469294 136294 469362 136350
rect 469418 136294 469488 136350
rect 469168 136226 469488 136294
rect 469168 136170 469238 136226
rect 469294 136170 469362 136226
rect 469418 136170 469488 136226
rect 469168 136102 469488 136170
rect 469168 136046 469238 136102
rect 469294 136046 469362 136102
rect 469418 136046 469488 136102
rect 469168 135978 469488 136046
rect 469168 135922 469238 135978
rect 469294 135922 469362 135978
rect 469418 135922 469488 135978
rect 469168 135888 469488 135922
rect 499888 136350 500208 136384
rect 499888 136294 499958 136350
rect 500014 136294 500082 136350
rect 500138 136294 500208 136350
rect 499888 136226 500208 136294
rect 499888 136170 499958 136226
rect 500014 136170 500082 136226
rect 500138 136170 500208 136226
rect 499888 136102 500208 136170
rect 499888 136046 499958 136102
rect 500014 136046 500082 136102
rect 500138 136046 500208 136102
rect 499888 135978 500208 136046
rect 499888 135922 499958 135978
rect 500014 135922 500082 135978
rect 500138 135922 500208 135978
rect 499888 135888 500208 135922
rect 530608 136350 530928 136384
rect 530608 136294 530678 136350
rect 530734 136294 530802 136350
rect 530858 136294 530928 136350
rect 530608 136226 530928 136294
rect 530608 136170 530678 136226
rect 530734 136170 530802 136226
rect 530858 136170 530928 136226
rect 530608 136102 530928 136170
rect 530608 136046 530678 136102
rect 530734 136046 530802 136102
rect 530858 136046 530928 136102
rect 530608 135978 530928 136046
rect 530608 135922 530678 135978
rect 530734 135922 530802 135978
rect 530858 135922 530928 135978
rect 530608 135888 530928 135922
rect 111154 130294 111250 130350
rect 111306 130294 111374 130350
rect 111430 130294 111498 130350
rect 111554 130294 111622 130350
rect 111678 130294 111774 130350
rect 111154 130226 111774 130294
rect 111154 130170 111250 130226
rect 111306 130170 111374 130226
rect 111430 130170 111498 130226
rect 111554 130170 111622 130226
rect 111678 130170 111774 130226
rect 111154 130102 111774 130170
rect 111154 130046 111250 130102
rect 111306 130046 111374 130102
rect 111430 130046 111498 130102
rect 111554 130046 111622 130102
rect 111678 130046 111774 130102
rect 111154 129978 111774 130046
rect 111154 129922 111250 129978
rect 111306 129922 111374 129978
rect 111430 129922 111498 129978
rect 111554 129922 111622 129978
rect 111678 129922 111774 129978
rect 96874 118294 96970 118350
rect 97026 118294 97094 118350
rect 97150 118294 97218 118350
rect 97274 118294 97342 118350
rect 97398 118294 97494 118350
rect 96874 118226 97494 118294
rect 96874 118170 96970 118226
rect 97026 118170 97094 118226
rect 97150 118170 97218 118226
rect 97274 118170 97342 118226
rect 97398 118170 97494 118226
rect 96874 118102 97494 118170
rect 96874 118046 96970 118102
rect 97026 118046 97094 118102
rect 97150 118046 97218 118102
rect 97274 118046 97342 118102
rect 97398 118046 97494 118102
rect 96874 117978 97494 118046
rect 96874 117922 96970 117978
rect 97026 117922 97094 117978
rect 97150 117922 97218 117978
rect 97274 117922 97342 117978
rect 97398 117922 97494 117978
rect 96874 100350 97494 117922
rect 100528 118350 100848 118384
rect 100528 118294 100598 118350
rect 100654 118294 100722 118350
rect 100778 118294 100848 118350
rect 100528 118226 100848 118294
rect 100528 118170 100598 118226
rect 100654 118170 100722 118226
rect 100778 118170 100848 118226
rect 100528 118102 100848 118170
rect 100528 118046 100598 118102
rect 100654 118046 100722 118102
rect 100778 118046 100848 118102
rect 100528 117978 100848 118046
rect 100528 117922 100598 117978
rect 100654 117922 100722 117978
rect 100778 117922 100848 117978
rect 100528 117888 100848 117922
rect 111154 112350 111774 129922
rect 115888 130350 116208 130384
rect 115888 130294 115958 130350
rect 116014 130294 116082 130350
rect 116138 130294 116208 130350
rect 115888 130226 116208 130294
rect 115888 130170 115958 130226
rect 116014 130170 116082 130226
rect 116138 130170 116208 130226
rect 115888 130102 116208 130170
rect 115888 130046 115958 130102
rect 116014 130046 116082 130102
rect 116138 130046 116208 130102
rect 115888 129978 116208 130046
rect 115888 129922 115958 129978
rect 116014 129922 116082 129978
rect 116138 129922 116208 129978
rect 115888 129888 116208 129922
rect 146608 130350 146928 130384
rect 146608 130294 146678 130350
rect 146734 130294 146802 130350
rect 146858 130294 146928 130350
rect 146608 130226 146928 130294
rect 146608 130170 146678 130226
rect 146734 130170 146802 130226
rect 146858 130170 146928 130226
rect 146608 130102 146928 130170
rect 146608 130046 146678 130102
rect 146734 130046 146802 130102
rect 146858 130046 146928 130102
rect 146608 129978 146928 130046
rect 146608 129922 146678 129978
rect 146734 129922 146802 129978
rect 146858 129922 146928 129978
rect 146608 129888 146928 129922
rect 177328 130350 177648 130384
rect 177328 130294 177398 130350
rect 177454 130294 177522 130350
rect 177578 130294 177648 130350
rect 177328 130226 177648 130294
rect 177328 130170 177398 130226
rect 177454 130170 177522 130226
rect 177578 130170 177648 130226
rect 177328 130102 177648 130170
rect 177328 130046 177398 130102
rect 177454 130046 177522 130102
rect 177578 130046 177648 130102
rect 177328 129978 177648 130046
rect 177328 129922 177398 129978
rect 177454 129922 177522 129978
rect 177578 129922 177648 129978
rect 177328 129888 177648 129922
rect 208048 130350 208368 130384
rect 208048 130294 208118 130350
rect 208174 130294 208242 130350
rect 208298 130294 208368 130350
rect 208048 130226 208368 130294
rect 208048 130170 208118 130226
rect 208174 130170 208242 130226
rect 208298 130170 208368 130226
rect 208048 130102 208368 130170
rect 208048 130046 208118 130102
rect 208174 130046 208242 130102
rect 208298 130046 208368 130102
rect 208048 129978 208368 130046
rect 208048 129922 208118 129978
rect 208174 129922 208242 129978
rect 208298 129922 208368 129978
rect 208048 129888 208368 129922
rect 238768 130350 239088 130384
rect 238768 130294 238838 130350
rect 238894 130294 238962 130350
rect 239018 130294 239088 130350
rect 238768 130226 239088 130294
rect 238768 130170 238838 130226
rect 238894 130170 238962 130226
rect 239018 130170 239088 130226
rect 238768 130102 239088 130170
rect 238768 130046 238838 130102
rect 238894 130046 238962 130102
rect 239018 130046 239088 130102
rect 238768 129978 239088 130046
rect 238768 129922 238838 129978
rect 238894 129922 238962 129978
rect 239018 129922 239088 129978
rect 238768 129888 239088 129922
rect 269488 130350 269808 130384
rect 269488 130294 269558 130350
rect 269614 130294 269682 130350
rect 269738 130294 269808 130350
rect 269488 130226 269808 130294
rect 269488 130170 269558 130226
rect 269614 130170 269682 130226
rect 269738 130170 269808 130226
rect 269488 130102 269808 130170
rect 269488 130046 269558 130102
rect 269614 130046 269682 130102
rect 269738 130046 269808 130102
rect 269488 129978 269808 130046
rect 269488 129922 269558 129978
rect 269614 129922 269682 129978
rect 269738 129922 269808 129978
rect 269488 129888 269808 129922
rect 300208 130350 300528 130384
rect 300208 130294 300278 130350
rect 300334 130294 300402 130350
rect 300458 130294 300528 130350
rect 300208 130226 300528 130294
rect 300208 130170 300278 130226
rect 300334 130170 300402 130226
rect 300458 130170 300528 130226
rect 300208 130102 300528 130170
rect 300208 130046 300278 130102
rect 300334 130046 300402 130102
rect 300458 130046 300528 130102
rect 300208 129978 300528 130046
rect 300208 129922 300278 129978
rect 300334 129922 300402 129978
rect 300458 129922 300528 129978
rect 300208 129888 300528 129922
rect 330928 130350 331248 130384
rect 330928 130294 330998 130350
rect 331054 130294 331122 130350
rect 331178 130294 331248 130350
rect 330928 130226 331248 130294
rect 330928 130170 330998 130226
rect 331054 130170 331122 130226
rect 331178 130170 331248 130226
rect 330928 130102 331248 130170
rect 330928 130046 330998 130102
rect 331054 130046 331122 130102
rect 331178 130046 331248 130102
rect 330928 129978 331248 130046
rect 330928 129922 330998 129978
rect 331054 129922 331122 129978
rect 331178 129922 331248 129978
rect 330928 129888 331248 129922
rect 361648 130350 361968 130384
rect 361648 130294 361718 130350
rect 361774 130294 361842 130350
rect 361898 130294 361968 130350
rect 361648 130226 361968 130294
rect 361648 130170 361718 130226
rect 361774 130170 361842 130226
rect 361898 130170 361968 130226
rect 361648 130102 361968 130170
rect 361648 130046 361718 130102
rect 361774 130046 361842 130102
rect 361898 130046 361968 130102
rect 361648 129978 361968 130046
rect 361648 129922 361718 129978
rect 361774 129922 361842 129978
rect 361898 129922 361968 129978
rect 361648 129888 361968 129922
rect 392368 130350 392688 130384
rect 392368 130294 392438 130350
rect 392494 130294 392562 130350
rect 392618 130294 392688 130350
rect 392368 130226 392688 130294
rect 392368 130170 392438 130226
rect 392494 130170 392562 130226
rect 392618 130170 392688 130226
rect 392368 130102 392688 130170
rect 392368 130046 392438 130102
rect 392494 130046 392562 130102
rect 392618 130046 392688 130102
rect 392368 129978 392688 130046
rect 392368 129922 392438 129978
rect 392494 129922 392562 129978
rect 392618 129922 392688 129978
rect 392368 129888 392688 129922
rect 423088 130350 423408 130384
rect 423088 130294 423158 130350
rect 423214 130294 423282 130350
rect 423338 130294 423408 130350
rect 423088 130226 423408 130294
rect 423088 130170 423158 130226
rect 423214 130170 423282 130226
rect 423338 130170 423408 130226
rect 423088 130102 423408 130170
rect 423088 130046 423158 130102
rect 423214 130046 423282 130102
rect 423338 130046 423408 130102
rect 423088 129978 423408 130046
rect 423088 129922 423158 129978
rect 423214 129922 423282 129978
rect 423338 129922 423408 129978
rect 423088 129888 423408 129922
rect 453808 130350 454128 130384
rect 453808 130294 453878 130350
rect 453934 130294 454002 130350
rect 454058 130294 454128 130350
rect 453808 130226 454128 130294
rect 453808 130170 453878 130226
rect 453934 130170 454002 130226
rect 454058 130170 454128 130226
rect 453808 130102 454128 130170
rect 453808 130046 453878 130102
rect 453934 130046 454002 130102
rect 454058 130046 454128 130102
rect 453808 129978 454128 130046
rect 453808 129922 453878 129978
rect 453934 129922 454002 129978
rect 454058 129922 454128 129978
rect 453808 129888 454128 129922
rect 484528 130350 484848 130384
rect 484528 130294 484598 130350
rect 484654 130294 484722 130350
rect 484778 130294 484848 130350
rect 484528 130226 484848 130294
rect 484528 130170 484598 130226
rect 484654 130170 484722 130226
rect 484778 130170 484848 130226
rect 484528 130102 484848 130170
rect 484528 130046 484598 130102
rect 484654 130046 484722 130102
rect 484778 130046 484848 130102
rect 484528 129978 484848 130046
rect 484528 129922 484598 129978
rect 484654 129922 484722 129978
rect 484778 129922 484848 129978
rect 484528 129888 484848 129922
rect 515248 130350 515568 130384
rect 515248 130294 515318 130350
rect 515374 130294 515442 130350
rect 515498 130294 515568 130350
rect 515248 130226 515568 130294
rect 515248 130170 515318 130226
rect 515374 130170 515442 130226
rect 515498 130170 515568 130226
rect 515248 130102 515568 130170
rect 515248 130046 515318 130102
rect 515374 130046 515442 130102
rect 515498 130046 515568 130102
rect 515248 129978 515568 130046
rect 515248 129922 515318 129978
rect 515374 129922 515442 129978
rect 515498 129922 515568 129978
rect 515248 129888 515568 129922
rect 545968 130350 546288 130384
rect 545968 130294 546038 130350
rect 546094 130294 546162 130350
rect 546218 130294 546288 130350
rect 545968 130226 546288 130294
rect 545968 130170 546038 130226
rect 546094 130170 546162 130226
rect 546218 130170 546288 130226
rect 545968 130102 546288 130170
rect 545968 130046 546038 130102
rect 546094 130046 546162 130102
rect 546218 130046 546288 130102
rect 545968 129978 546288 130046
rect 545968 129922 546038 129978
rect 546094 129922 546162 129978
rect 546218 129922 546288 129978
rect 545968 129888 546288 129922
rect 561154 130350 561774 147922
rect 561154 130294 561250 130350
rect 561306 130294 561374 130350
rect 561430 130294 561498 130350
rect 561554 130294 561622 130350
rect 561678 130294 561774 130350
rect 561154 130226 561774 130294
rect 561154 130170 561250 130226
rect 561306 130170 561374 130226
rect 561430 130170 561498 130226
rect 561554 130170 561622 130226
rect 561678 130170 561774 130226
rect 561154 130102 561774 130170
rect 561154 130046 561250 130102
rect 561306 130046 561374 130102
rect 561430 130046 561498 130102
rect 561554 130046 561622 130102
rect 561678 130046 561774 130102
rect 561154 129978 561774 130046
rect 561154 129922 561250 129978
rect 561306 129922 561374 129978
rect 561430 129922 561498 129978
rect 561554 129922 561622 129978
rect 561678 129922 561774 129978
rect 131248 118350 131568 118384
rect 131248 118294 131318 118350
rect 131374 118294 131442 118350
rect 131498 118294 131568 118350
rect 131248 118226 131568 118294
rect 131248 118170 131318 118226
rect 131374 118170 131442 118226
rect 131498 118170 131568 118226
rect 131248 118102 131568 118170
rect 131248 118046 131318 118102
rect 131374 118046 131442 118102
rect 131498 118046 131568 118102
rect 131248 117978 131568 118046
rect 131248 117922 131318 117978
rect 131374 117922 131442 117978
rect 131498 117922 131568 117978
rect 131248 117888 131568 117922
rect 161968 118350 162288 118384
rect 161968 118294 162038 118350
rect 162094 118294 162162 118350
rect 162218 118294 162288 118350
rect 161968 118226 162288 118294
rect 161968 118170 162038 118226
rect 162094 118170 162162 118226
rect 162218 118170 162288 118226
rect 161968 118102 162288 118170
rect 161968 118046 162038 118102
rect 162094 118046 162162 118102
rect 162218 118046 162288 118102
rect 161968 117978 162288 118046
rect 161968 117922 162038 117978
rect 162094 117922 162162 117978
rect 162218 117922 162288 117978
rect 161968 117888 162288 117922
rect 192688 118350 193008 118384
rect 192688 118294 192758 118350
rect 192814 118294 192882 118350
rect 192938 118294 193008 118350
rect 192688 118226 193008 118294
rect 192688 118170 192758 118226
rect 192814 118170 192882 118226
rect 192938 118170 193008 118226
rect 192688 118102 193008 118170
rect 192688 118046 192758 118102
rect 192814 118046 192882 118102
rect 192938 118046 193008 118102
rect 192688 117978 193008 118046
rect 192688 117922 192758 117978
rect 192814 117922 192882 117978
rect 192938 117922 193008 117978
rect 192688 117888 193008 117922
rect 223408 118350 223728 118384
rect 223408 118294 223478 118350
rect 223534 118294 223602 118350
rect 223658 118294 223728 118350
rect 223408 118226 223728 118294
rect 223408 118170 223478 118226
rect 223534 118170 223602 118226
rect 223658 118170 223728 118226
rect 223408 118102 223728 118170
rect 223408 118046 223478 118102
rect 223534 118046 223602 118102
rect 223658 118046 223728 118102
rect 223408 117978 223728 118046
rect 223408 117922 223478 117978
rect 223534 117922 223602 117978
rect 223658 117922 223728 117978
rect 223408 117888 223728 117922
rect 254128 118350 254448 118384
rect 254128 118294 254198 118350
rect 254254 118294 254322 118350
rect 254378 118294 254448 118350
rect 254128 118226 254448 118294
rect 254128 118170 254198 118226
rect 254254 118170 254322 118226
rect 254378 118170 254448 118226
rect 254128 118102 254448 118170
rect 254128 118046 254198 118102
rect 254254 118046 254322 118102
rect 254378 118046 254448 118102
rect 254128 117978 254448 118046
rect 254128 117922 254198 117978
rect 254254 117922 254322 117978
rect 254378 117922 254448 117978
rect 254128 117888 254448 117922
rect 284848 118350 285168 118384
rect 284848 118294 284918 118350
rect 284974 118294 285042 118350
rect 285098 118294 285168 118350
rect 284848 118226 285168 118294
rect 284848 118170 284918 118226
rect 284974 118170 285042 118226
rect 285098 118170 285168 118226
rect 284848 118102 285168 118170
rect 284848 118046 284918 118102
rect 284974 118046 285042 118102
rect 285098 118046 285168 118102
rect 284848 117978 285168 118046
rect 284848 117922 284918 117978
rect 284974 117922 285042 117978
rect 285098 117922 285168 117978
rect 284848 117888 285168 117922
rect 315568 118350 315888 118384
rect 315568 118294 315638 118350
rect 315694 118294 315762 118350
rect 315818 118294 315888 118350
rect 315568 118226 315888 118294
rect 315568 118170 315638 118226
rect 315694 118170 315762 118226
rect 315818 118170 315888 118226
rect 315568 118102 315888 118170
rect 315568 118046 315638 118102
rect 315694 118046 315762 118102
rect 315818 118046 315888 118102
rect 315568 117978 315888 118046
rect 315568 117922 315638 117978
rect 315694 117922 315762 117978
rect 315818 117922 315888 117978
rect 315568 117888 315888 117922
rect 346288 118350 346608 118384
rect 346288 118294 346358 118350
rect 346414 118294 346482 118350
rect 346538 118294 346608 118350
rect 346288 118226 346608 118294
rect 346288 118170 346358 118226
rect 346414 118170 346482 118226
rect 346538 118170 346608 118226
rect 346288 118102 346608 118170
rect 346288 118046 346358 118102
rect 346414 118046 346482 118102
rect 346538 118046 346608 118102
rect 346288 117978 346608 118046
rect 346288 117922 346358 117978
rect 346414 117922 346482 117978
rect 346538 117922 346608 117978
rect 346288 117888 346608 117922
rect 377008 118350 377328 118384
rect 377008 118294 377078 118350
rect 377134 118294 377202 118350
rect 377258 118294 377328 118350
rect 377008 118226 377328 118294
rect 377008 118170 377078 118226
rect 377134 118170 377202 118226
rect 377258 118170 377328 118226
rect 377008 118102 377328 118170
rect 377008 118046 377078 118102
rect 377134 118046 377202 118102
rect 377258 118046 377328 118102
rect 377008 117978 377328 118046
rect 377008 117922 377078 117978
rect 377134 117922 377202 117978
rect 377258 117922 377328 117978
rect 377008 117888 377328 117922
rect 407728 118350 408048 118384
rect 407728 118294 407798 118350
rect 407854 118294 407922 118350
rect 407978 118294 408048 118350
rect 407728 118226 408048 118294
rect 407728 118170 407798 118226
rect 407854 118170 407922 118226
rect 407978 118170 408048 118226
rect 407728 118102 408048 118170
rect 407728 118046 407798 118102
rect 407854 118046 407922 118102
rect 407978 118046 408048 118102
rect 407728 117978 408048 118046
rect 407728 117922 407798 117978
rect 407854 117922 407922 117978
rect 407978 117922 408048 117978
rect 407728 117888 408048 117922
rect 438448 118350 438768 118384
rect 438448 118294 438518 118350
rect 438574 118294 438642 118350
rect 438698 118294 438768 118350
rect 438448 118226 438768 118294
rect 438448 118170 438518 118226
rect 438574 118170 438642 118226
rect 438698 118170 438768 118226
rect 438448 118102 438768 118170
rect 438448 118046 438518 118102
rect 438574 118046 438642 118102
rect 438698 118046 438768 118102
rect 438448 117978 438768 118046
rect 438448 117922 438518 117978
rect 438574 117922 438642 117978
rect 438698 117922 438768 117978
rect 438448 117888 438768 117922
rect 469168 118350 469488 118384
rect 469168 118294 469238 118350
rect 469294 118294 469362 118350
rect 469418 118294 469488 118350
rect 469168 118226 469488 118294
rect 469168 118170 469238 118226
rect 469294 118170 469362 118226
rect 469418 118170 469488 118226
rect 469168 118102 469488 118170
rect 469168 118046 469238 118102
rect 469294 118046 469362 118102
rect 469418 118046 469488 118102
rect 469168 117978 469488 118046
rect 469168 117922 469238 117978
rect 469294 117922 469362 117978
rect 469418 117922 469488 117978
rect 469168 117888 469488 117922
rect 499888 118350 500208 118384
rect 499888 118294 499958 118350
rect 500014 118294 500082 118350
rect 500138 118294 500208 118350
rect 499888 118226 500208 118294
rect 499888 118170 499958 118226
rect 500014 118170 500082 118226
rect 500138 118170 500208 118226
rect 499888 118102 500208 118170
rect 499888 118046 499958 118102
rect 500014 118046 500082 118102
rect 500138 118046 500208 118102
rect 499888 117978 500208 118046
rect 499888 117922 499958 117978
rect 500014 117922 500082 117978
rect 500138 117922 500208 117978
rect 499888 117888 500208 117922
rect 530608 118350 530928 118384
rect 530608 118294 530678 118350
rect 530734 118294 530802 118350
rect 530858 118294 530928 118350
rect 530608 118226 530928 118294
rect 530608 118170 530678 118226
rect 530734 118170 530802 118226
rect 530858 118170 530928 118226
rect 530608 118102 530928 118170
rect 530608 118046 530678 118102
rect 530734 118046 530802 118102
rect 530858 118046 530928 118102
rect 530608 117978 530928 118046
rect 530608 117922 530678 117978
rect 530734 117922 530802 117978
rect 530858 117922 530928 117978
rect 530608 117888 530928 117922
rect 111154 112294 111250 112350
rect 111306 112294 111374 112350
rect 111430 112294 111498 112350
rect 111554 112294 111622 112350
rect 111678 112294 111774 112350
rect 111154 112226 111774 112294
rect 111154 112170 111250 112226
rect 111306 112170 111374 112226
rect 111430 112170 111498 112226
rect 111554 112170 111622 112226
rect 111678 112170 111774 112226
rect 111154 112102 111774 112170
rect 111154 112046 111250 112102
rect 111306 112046 111374 112102
rect 111430 112046 111498 112102
rect 111554 112046 111622 112102
rect 111678 112046 111774 112102
rect 111154 111978 111774 112046
rect 111154 111922 111250 111978
rect 111306 111922 111374 111978
rect 111430 111922 111498 111978
rect 111554 111922 111622 111978
rect 111678 111922 111774 111978
rect 96874 100294 96970 100350
rect 97026 100294 97094 100350
rect 97150 100294 97218 100350
rect 97274 100294 97342 100350
rect 97398 100294 97494 100350
rect 96874 100226 97494 100294
rect 96874 100170 96970 100226
rect 97026 100170 97094 100226
rect 97150 100170 97218 100226
rect 97274 100170 97342 100226
rect 97398 100170 97494 100226
rect 96874 100102 97494 100170
rect 96874 100046 96970 100102
rect 97026 100046 97094 100102
rect 97150 100046 97218 100102
rect 97274 100046 97342 100102
rect 97398 100046 97494 100102
rect 96874 99978 97494 100046
rect 96874 99922 96970 99978
rect 97026 99922 97094 99978
rect 97150 99922 97218 99978
rect 97274 99922 97342 99978
rect 97398 99922 97494 99978
rect 96874 82350 97494 99922
rect 100528 100350 100848 100384
rect 100528 100294 100598 100350
rect 100654 100294 100722 100350
rect 100778 100294 100848 100350
rect 100528 100226 100848 100294
rect 100528 100170 100598 100226
rect 100654 100170 100722 100226
rect 100778 100170 100848 100226
rect 100528 100102 100848 100170
rect 100528 100046 100598 100102
rect 100654 100046 100722 100102
rect 100778 100046 100848 100102
rect 100528 99978 100848 100046
rect 100528 99922 100598 99978
rect 100654 99922 100722 99978
rect 100778 99922 100848 99978
rect 100528 99888 100848 99922
rect 111154 94350 111774 111922
rect 115888 112350 116208 112384
rect 115888 112294 115958 112350
rect 116014 112294 116082 112350
rect 116138 112294 116208 112350
rect 115888 112226 116208 112294
rect 115888 112170 115958 112226
rect 116014 112170 116082 112226
rect 116138 112170 116208 112226
rect 115888 112102 116208 112170
rect 115888 112046 115958 112102
rect 116014 112046 116082 112102
rect 116138 112046 116208 112102
rect 115888 111978 116208 112046
rect 115888 111922 115958 111978
rect 116014 111922 116082 111978
rect 116138 111922 116208 111978
rect 115888 111888 116208 111922
rect 146608 112350 146928 112384
rect 146608 112294 146678 112350
rect 146734 112294 146802 112350
rect 146858 112294 146928 112350
rect 146608 112226 146928 112294
rect 146608 112170 146678 112226
rect 146734 112170 146802 112226
rect 146858 112170 146928 112226
rect 146608 112102 146928 112170
rect 146608 112046 146678 112102
rect 146734 112046 146802 112102
rect 146858 112046 146928 112102
rect 146608 111978 146928 112046
rect 146608 111922 146678 111978
rect 146734 111922 146802 111978
rect 146858 111922 146928 111978
rect 146608 111888 146928 111922
rect 177328 112350 177648 112384
rect 177328 112294 177398 112350
rect 177454 112294 177522 112350
rect 177578 112294 177648 112350
rect 177328 112226 177648 112294
rect 177328 112170 177398 112226
rect 177454 112170 177522 112226
rect 177578 112170 177648 112226
rect 177328 112102 177648 112170
rect 177328 112046 177398 112102
rect 177454 112046 177522 112102
rect 177578 112046 177648 112102
rect 177328 111978 177648 112046
rect 177328 111922 177398 111978
rect 177454 111922 177522 111978
rect 177578 111922 177648 111978
rect 177328 111888 177648 111922
rect 208048 112350 208368 112384
rect 208048 112294 208118 112350
rect 208174 112294 208242 112350
rect 208298 112294 208368 112350
rect 208048 112226 208368 112294
rect 208048 112170 208118 112226
rect 208174 112170 208242 112226
rect 208298 112170 208368 112226
rect 208048 112102 208368 112170
rect 208048 112046 208118 112102
rect 208174 112046 208242 112102
rect 208298 112046 208368 112102
rect 208048 111978 208368 112046
rect 208048 111922 208118 111978
rect 208174 111922 208242 111978
rect 208298 111922 208368 111978
rect 208048 111888 208368 111922
rect 238768 112350 239088 112384
rect 238768 112294 238838 112350
rect 238894 112294 238962 112350
rect 239018 112294 239088 112350
rect 238768 112226 239088 112294
rect 238768 112170 238838 112226
rect 238894 112170 238962 112226
rect 239018 112170 239088 112226
rect 238768 112102 239088 112170
rect 238768 112046 238838 112102
rect 238894 112046 238962 112102
rect 239018 112046 239088 112102
rect 238768 111978 239088 112046
rect 238768 111922 238838 111978
rect 238894 111922 238962 111978
rect 239018 111922 239088 111978
rect 238768 111888 239088 111922
rect 269488 112350 269808 112384
rect 269488 112294 269558 112350
rect 269614 112294 269682 112350
rect 269738 112294 269808 112350
rect 269488 112226 269808 112294
rect 269488 112170 269558 112226
rect 269614 112170 269682 112226
rect 269738 112170 269808 112226
rect 269488 112102 269808 112170
rect 269488 112046 269558 112102
rect 269614 112046 269682 112102
rect 269738 112046 269808 112102
rect 269488 111978 269808 112046
rect 269488 111922 269558 111978
rect 269614 111922 269682 111978
rect 269738 111922 269808 111978
rect 269488 111888 269808 111922
rect 300208 112350 300528 112384
rect 300208 112294 300278 112350
rect 300334 112294 300402 112350
rect 300458 112294 300528 112350
rect 300208 112226 300528 112294
rect 300208 112170 300278 112226
rect 300334 112170 300402 112226
rect 300458 112170 300528 112226
rect 300208 112102 300528 112170
rect 300208 112046 300278 112102
rect 300334 112046 300402 112102
rect 300458 112046 300528 112102
rect 300208 111978 300528 112046
rect 300208 111922 300278 111978
rect 300334 111922 300402 111978
rect 300458 111922 300528 111978
rect 300208 111888 300528 111922
rect 330928 112350 331248 112384
rect 330928 112294 330998 112350
rect 331054 112294 331122 112350
rect 331178 112294 331248 112350
rect 330928 112226 331248 112294
rect 330928 112170 330998 112226
rect 331054 112170 331122 112226
rect 331178 112170 331248 112226
rect 330928 112102 331248 112170
rect 330928 112046 330998 112102
rect 331054 112046 331122 112102
rect 331178 112046 331248 112102
rect 330928 111978 331248 112046
rect 330928 111922 330998 111978
rect 331054 111922 331122 111978
rect 331178 111922 331248 111978
rect 330928 111888 331248 111922
rect 361648 112350 361968 112384
rect 361648 112294 361718 112350
rect 361774 112294 361842 112350
rect 361898 112294 361968 112350
rect 361648 112226 361968 112294
rect 361648 112170 361718 112226
rect 361774 112170 361842 112226
rect 361898 112170 361968 112226
rect 361648 112102 361968 112170
rect 361648 112046 361718 112102
rect 361774 112046 361842 112102
rect 361898 112046 361968 112102
rect 361648 111978 361968 112046
rect 361648 111922 361718 111978
rect 361774 111922 361842 111978
rect 361898 111922 361968 111978
rect 361648 111888 361968 111922
rect 392368 112350 392688 112384
rect 392368 112294 392438 112350
rect 392494 112294 392562 112350
rect 392618 112294 392688 112350
rect 392368 112226 392688 112294
rect 392368 112170 392438 112226
rect 392494 112170 392562 112226
rect 392618 112170 392688 112226
rect 392368 112102 392688 112170
rect 392368 112046 392438 112102
rect 392494 112046 392562 112102
rect 392618 112046 392688 112102
rect 392368 111978 392688 112046
rect 392368 111922 392438 111978
rect 392494 111922 392562 111978
rect 392618 111922 392688 111978
rect 392368 111888 392688 111922
rect 423088 112350 423408 112384
rect 423088 112294 423158 112350
rect 423214 112294 423282 112350
rect 423338 112294 423408 112350
rect 423088 112226 423408 112294
rect 423088 112170 423158 112226
rect 423214 112170 423282 112226
rect 423338 112170 423408 112226
rect 423088 112102 423408 112170
rect 423088 112046 423158 112102
rect 423214 112046 423282 112102
rect 423338 112046 423408 112102
rect 423088 111978 423408 112046
rect 423088 111922 423158 111978
rect 423214 111922 423282 111978
rect 423338 111922 423408 111978
rect 423088 111888 423408 111922
rect 453808 112350 454128 112384
rect 453808 112294 453878 112350
rect 453934 112294 454002 112350
rect 454058 112294 454128 112350
rect 453808 112226 454128 112294
rect 453808 112170 453878 112226
rect 453934 112170 454002 112226
rect 454058 112170 454128 112226
rect 453808 112102 454128 112170
rect 453808 112046 453878 112102
rect 453934 112046 454002 112102
rect 454058 112046 454128 112102
rect 453808 111978 454128 112046
rect 453808 111922 453878 111978
rect 453934 111922 454002 111978
rect 454058 111922 454128 111978
rect 453808 111888 454128 111922
rect 484528 112350 484848 112384
rect 484528 112294 484598 112350
rect 484654 112294 484722 112350
rect 484778 112294 484848 112350
rect 484528 112226 484848 112294
rect 484528 112170 484598 112226
rect 484654 112170 484722 112226
rect 484778 112170 484848 112226
rect 484528 112102 484848 112170
rect 484528 112046 484598 112102
rect 484654 112046 484722 112102
rect 484778 112046 484848 112102
rect 484528 111978 484848 112046
rect 484528 111922 484598 111978
rect 484654 111922 484722 111978
rect 484778 111922 484848 111978
rect 484528 111888 484848 111922
rect 515248 112350 515568 112384
rect 515248 112294 515318 112350
rect 515374 112294 515442 112350
rect 515498 112294 515568 112350
rect 515248 112226 515568 112294
rect 515248 112170 515318 112226
rect 515374 112170 515442 112226
rect 515498 112170 515568 112226
rect 515248 112102 515568 112170
rect 515248 112046 515318 112102
rect 515374 112046 515442 112102
rect 515498 112046 515568 112102
rect 515248 111978 515568 112046
rect 515248 111922 515318 111978
rect 515374 111922 515442 111978
rect 515498 111922 515568 111978
rect 515248 111888 515568 111922
rect 545968 112350 546288 112384
rect 545968 112294 546038 112350
rect 546094 112294 546162 112350
rect 546218 112294 546288 112350
rect 545968 112226 546288 112294
rect 545968 112170 546038 112226
rect 546094 112170 546162 112226
rect 546218 112170 546288 112226
rect 545968 112102 546288 112170
rect 545968 112046 546038 112102
rect 546094 112046 546162 112102
rect 546218 112046 546288 112102
rect 545968 111978 546288 112046
rect 545968 111922 546038 111978
rect 546094 111922 546162 111978
rect 546218 111922 546288 111978
rect 545968 111888 546288 111922
rect 561154 112350 561774 129922
rect 561154 112294 561250 112350
rect 561306 112294 561374 112350
rect 561430 112294 561498 112350
rect 561554 112294 561622 112350
rect 561678 112294 561774 112350
rect 561154 112226 561774 112294
rect 561154 112170 561250 112226
rect 561306 112170 561374 112226
rect 561430 112170 561498 112226
rect 561554 112170 561622 112226
rect 561678 112170 561774 112226
rect 561154 112102 561774 112170
rect 561154 112046 561250 112102
rect 561306 112046 561374 112102
rect 561430 112046 561498 112102
rect 561554 112046 561622 112102
rect 561678 112046 561774 112102
rect 561154 111978 561774 112046
rect 561154 111922 561250 111978
rect 561306 111922 561374 111978
rect 561430 111922 561498 111978
rect 561554 111922 561622 111978
rect 561678 111922 561774 111978
rect 131248 100350 131568 100384
rect 131248 100294 131318 100350
rect 131374 100294 131442 100350
rect 131498 100294 131568 100350
rect 131248 100226 131568 100294
rect 131248 100170 131318 100226
rect 131374 100170 131442 100226
rect 131498 100170 131568 100226
rect 131248 100102 131568 100170
rect 131248 100046 131318 100102
rect 131374 100046 131442 100102
rect 131498 100046 131568 100102
rect 131248 99978 131568 100046
rect 131248 99922 131318 99978
rect 131374 99922 131442 99978
rect 131498 99922 131568 99978
rect 131248 99888 131568 99922
rect 161968 100350 162288 100384
rect 161968 100294 162038 100350
rect 162094 100294 162162 100350
rect 162218 100294 162288 100350
rect 161968 100226 162288 100294
rect 161968 100170 162038 100226
rect 162094 100170 162162 100226
rect 162218 100170 162288 100226
rect 161968 100102 162288 100170
rect 161968 100046 162038 100102
rect 162094 100046 162162 100102
rect 162218 100046 162288 100102
rect 161968 99978 162288 100046
rect 161968 99922 162038 99978
rect 162094 99922 162162 99978
rect 162218 99922 162288 99978
rect 161968 99888 162288 99922
rect 192688 100350 193008 100384
rect 192688 100294 192758 100350
rect 192814 100294 192882 100350
rect 192938 100294 193008 100350
rect 192688 100226 193008 100294
rect 192688 100170 192758 100226
rect 192814 100170 192882 100226
rect 192938 100170 193008 100226
rect 192688 100102 193008 100170
rect 192688 100046 192758 100102
rect 192814 100046 192882 100102
rect 192938 100046 193008 100102
rect 192688 99978 193008 100046
rect 192688 99922 192758 99978
rect 192814 99922 192882 99978
rect 192938 99922 193008 99978
rect 192688 99888 193008 99922
rect 223408 100350 223728 100384
rect 223408 100294 223478 100350
rect 223534 100294 223602 100350
rect 223658 100294 223728 100350
rect 223408 100226 223728 100294
rect 223408 100170 223478 100226
rect 223534 100170 223602 100226
rect 223658 100170 223728 100226
rect 223408 100102 223728 100170
rect 223408 100046 223478 100102
rect 223534 100046 223602 100102
rect 223658 100046 223728 100102
rect 223408 99978 223728 100046
rect 223408 99922 223478 99978
rect 223534 99922 223602 99978
rect 223658 99922 223728 99978
rect 223408 99888 223728 99922
rect 254128 100350 254448 100384
rect 254128 100294 254198 100350
rect 254254 100294 254322 100350
rect 254378 100294 254448 100350
rect 254128 100226 254448 100294
rect 254128 100170 254198 100226
rect 254254 100170 254322 100226
rect 254378 100170 254448 100226
rect 254128 100102 254448 100170
rect 254128 100046 254198 100102
rect 254254 100046 254322 100102
rect 254378 100046 254448 100102
rect 254128 99978 254448 100046
rect 254128 99922 254198 99978
rect 254254 99922 254322 99978
rect 254378 99922 254448 99978
rect 254128 99888 254448 99922
rect 284848 100350 285168 100384
rect 284848 100294 284918 100350
rect 284974 100294 285042 100350
rect 285098 100294 285168 100350
rect 284848 100226 285168 100294
rect 284848 100170 284918 100226
rect 284974 100170 285042 100226
rect 285098 100170 285168 100226
rect 284848 100102 285168 100170
rect 284848 100046 284918 100102
rect 284974 100046 285042 100102
rect 285098 100046 285168 100102
rect 284848 99978 285168 100046
rect 284848 99922 284918 99978
rect 284974 99922 285042 99978
rect 285098 99922 285168 99978
rect 284848 99888 285168 99922
rect 315568 100350 315888 100384
rect 315568 100294 315638 100350
rect 315694 100294 315762 100350
rect 315818 100294 315888 100350
rect 315568 100226 315888 100294
rect 315568 100170 315638 100226
rect 315694 100170 315762 100226
rect 315818 100170 315888 100226
rect 315568 100102 315888 100170
rect 315568 100046 315638 100102
rect 315694 100046 315762 100102
rect 315818 100046 315888 100102
rect 315568 99978 315888 100046
rect 315568 99922 315638 99978
rect 315694 99922 315762 99978
rect 315818 99922 315888 99978
rect 315568 99888 315888 99922
rect 346288 100350 346608 100384
rect 346288 100294 346358 100350
rect 346414 100294 346482 100350
rect 346538 100294 346608 100350
rect 346288 100226 346608 100294
rect 346288 100170 346358 100226
rect 346414 100170 346482 100226
rect 346538 100170 346608 100226
rect 346288 100102 346608 100170
rect 346288 100046 346358 100102
rect 346414 100046 346482 100102
rect 346538 100046 346608 100102
rect 346288 99978 346608 100046
rect 346288 99922 346358 99978
rect 346414 99922 346482 99978
rect 346538 99922 346608 99978
rect 346288 99888 346608 99922
rect 377008 100350 377328 100384
rect 377008 100294 377078 100350
rect 377134 100294 377202 100350
rect 377258 100294 377328 100350
rect 377008 100226 377328 100294
rect 377008 100170 377078 100226
rect 377134 100170 377202 100226
rect 377258 100170 377328 100226
rect 377008 100102 377328 100170
rect 377008 100046 377078 100102
rect 377134 100046 377202 100102
rect 377258 100046 377328 100102
rect 377008 99978 377328 100046
rect 377008 99922 377078 99978
rect 377134 99922 377202 99978
rect 377258 99922 377328 99978
rect 377008 99888 377328 99922
rect 407728 100350 408048 100384
rect 407728 100294 407798 100350
rect 407854 100294 407922 100350
rect 407978 100294 408048 100350
rect 407728 100226 408048 100294
rect 407728 100170 407798 100226
rect 407854 100170 407922 100226
rect 407978 100170 408048 100226
rect 407728 100102 408048 100170
rect 407728 100046 407798 100102
rect 407854 100046 407922 100102
rect 407978 100046 408048 100102
rect 407728 99978 408048 100046
rect 407728 99922 407798 99978
rect 407854 99922 407922 99978
rect 407978 99922 408048 99978
rect 407728 99888 408048 99922
rect 438448 100350 438768 100384
rect 438448 100294 438518 100350
rect 438574 100294 438642 100350
rect 438698 100294 438768 100350
rect 438448 100226 438768 100294
rect 438448 100170 438518 100226
rect 438574 100170 438642 100226
rect 438698 100170 438768 100226
rect 438448 100102 438768 100170
rect 438448 100046 438518 100102
rect 438574 100046 438642 100102
rect 438698 100046 438768 100102
rect 438448 99978 438768 100046
rect 438448 99922 438518 99978
rect 438574 99922 438642 99978
rect 438698 99922 438768 99978
rect 438448 99888 438768 99922
rect 469168 100350 469488 100384
rect 469168 100294 469238 100350
rect 469294 100294 469362 100350
rect 469418 100294 469488 100350
rect 469168 100226 469488 100294
rect 469168 100170 469238 100226
rect 469294 100170 469362 100226
rect 469418 100170 469488 100226
rect 469168 100102 469488 100170
rect 469168 100046 469238 100102
rect 469294 100046 469362 100102
rect 469418 100046 469488 100102
rect 469168 99978 469488 100046
rect 469168 99922 469238 99978
rect 469294 99922 469362 99978
rect 469418 99922 469488 99978
rect 469168 99888 469488 99922
rect 499888 100350 500208 100384
rect 499888 100294 499958 100350
rect 500014 100294 500082 100350
rect 500138 100294 500208 100350
rect 499888 100226 500208 100294
rect 499888 100170 499958 100226
rect 500014 100170 500082 100226
rect 500138 100170 500208 100226
rect 499888 100102 500208 100170
rect 499888 100046 499958 100102
rect 500014 100046 500082 100102
rect 500138 100046 500208 100102
rect 499888 99978 500208 100046
rect 499888 99922 499958 99978
rect 500014 99922 500082 99978
rect 500138 99922 500208 99978
rect 499888 99888 500208 99922
rect 530608 100350 530928 100384
rect 530608 100294 530678 100350
rect 530734 100294 530802 100350
rect 530858 100294 530928 100350
rect 530608 100226 530928 100294
rect 530608 100170 530678 100226
rect 530734 100170 530802 100226
rect 530858 100170 530928 100226
rect 530608 100102 530928 100170
rect 530608 100046 530678 100102
rect 530734 100046 530802 100102
rect 530858 100046 530928 100102
rect 530608 99978 530928 100046
rect 530608 99922 530678 99978
rect 530734 99922 530802 99978
rect 530858 99922 530928 99978
rect 530608 99888 530928 99922
rect 111154 94294 111250 94350
rect 111306 94294 111374 94350
rect 111430 94294 111498 94350
rect 111554 94294 111622 94350
rect 111678 94294 111774 94350
rect 111154 94226 111774 94294
rect 111154 94170 111250 94226
rect 111306 94170 111374 94226
rect 111430 94170 111498 94226
rect 111554 94170 111622 94226
rect 111678 94170 111774 94226
rect 111154 94102 111774 94170
rect 111154 94046 111250 94102
rect 111306 94046 111374 94102
rect 111430 94046 111498 94102
rect 111554 94046 111622 94102
rect 111678 94046 111774 94102
rect 111154 93978 111774 94046
rect 111154 93922 111250 93978
rect 111306 93922 111374 93978
rect 111430 93922 111498 93978
rect 111554 93922 111622 93978
rect 111678 93922 111774 93978
rect 96874 82294 96970 82350
rect 97026 82294 97094 82350
rect 97150 82294 97218 82350
rect 97274 82294 97342 82350
rect 97398 82294 97494 82350
rect 96874 82226 97494 82294
rect 96874 82170 96970 82226
rect 97026 82170 97094 82226
rect 97150 82170 97218 82226
rect 97274 82170 97342 82226
rect 97398 82170 97494 82226
rect 96874 82102 97494 82170
rect 96874 82046 96970 82102
rect 97026 82046 97094 82102
rect 97150 82046 97218 82102
rect 97274 82046 97342 82102
rect 97398 82046 97494 82102
rect 96874 81978 97494 82046
rect 96874 81922 96970 81978
rect 97026 81922 97094 81978
rect 97150 81922 97218 81978
rect 97274 81922 97342 81978
rect 97398 81922 97494 81978
rect 96874 64350 97494 81922
rect 100528 82350 100848 82384
rect 100528 82294 100598 82350
rect 100654 82294 100722 82350
rect 100778 82294 100848 82350
rect 100528 82226 100848 82294
rect 100528 82170 100598 82226
rect 100654 82170 100722 82226
rect 100778 82170 100848 82226
rect 100528 82102 100848 82170
rect 100528 82046 100598 82102
rect 100654 82046 100722 82102
rect 100778 82046 100848 82102
rect 100528 81978 100848 82046
rect 100528 81922 100598 81978
rect 100654 81922 100722 81978
rect 100778 81922 100848 81978
rect 100528 81888 100848 81922
rect 111154 76350 111774 93922
rect 115888 94350 116208 94384
rect 115888 94294 115958 94350
rect 116014 94294 116082 94350
rect 116138 94294 116208 94350
rect 115888 94226 116208 94294
rect 115888 94170 115958 94226
rect 116014 94170 116082 94226
rect 116138 94170 116208 94226
rect 115888 94102 116208 94170
rect 115888 94046 115958 94102
rect 116014 94046 116082 94102
rect 116138 94046 116208 94102
rect 115888 93978 116208 94046
rect 115888 93922 115958 93978
rect 116014 93922 116082 93978
rect 116138 93922 116208 93978
rect 115888 93888 116208 93922
rect 146608 94350 146928 94384
rect 146608 94294 146678 94350
rect 146734 94294 146802 94350
rect 146858 94294 146928 94350
rect 146608 94226 146928 94294
rect 146608 94170 146678 94226
rect 146734 94170 146802 94226
rect 146858 94170 146928 94226
rect 146608 94102 146928 94170
rect 146608 94046 146678 94102
rect 146734 94046 146802 94102
rect 146858 94046 146928 94102
rect 146608 93978 146928 94046
rect 146608 93922 146678 93978
rect 146734 93922 146802 93978
rect 146858 93922 146928 93978
rect 146608 93888 146928 93922
rect 177328 94350 177648 94384
rect 177328 94294 177398 94350
rect 177454 94294 177522 94350
rect 177578 94294 177648 94350
rect 177328 94226 177648 94294
rect 177328 94170 177398 94226
rect 177454 94170 177522 94226
rect 177578 94170 177648 94226
rect 177328 94102 177648 94170
rect 177328 94046 177398 94102
rect 177454 94046 177522 94102
rect 177578 94046 177648 94102
rect 177328 93978 177648 94046
rect 177328 93922 177398 93978
rect 177454 93922 177522 93978
rect 177578 93922 177648 93978
rect 177328 93888 177648 93922
rect 208048 94350 208368 94384
rect 208048 94294 208118 94350
rect 208174 94294 208242 94350
rect 208298 94294 208368 94350
rect 208048 94226 208368 94294
rect 208048 94170 208118 94226
rect 208174 94170 208242 94226
rect 208298 94170 208368 94226
rect 208048 94102 208368 94170
rect 208048 94046 208118 94102
rect 208174 94046 208242 94102
rect 208298 94046 208368 94102
rect 208048 93978 208368 94046
rect 208048 93922 208118 93978
rect 208174 93922 208242 93978
rect 208298 93922 208368 93978
rect 208048 93888 208368 93922
rect 238768 94350 239088 94384
rect 238768 94294 238838 94350
rect 238894 94294 238962 94350
rect 239018 94294 239088 94350
rect 238768 94226 239088 94294
rect 238768 94170 238838 94226
rect 238894 94170 238962 94226
rect 239018 94170 239088 94226
rect 238768 94102 239088 94170
rect 238768 94046 238838 94102
rect 238894 94046 238962 94102
rect 239018 94046 239088 94102
rect 238768 93978 239088 94046
rect 238768 93922 238838 93978
rect 238894 93922 238962 93978
rect 239018 93922 239088 93978
rect 238768 93888 239088 93922
rect 269488 94350 269808 94384
rect 269488 94294 269558 94350
rect 269614 94294 269682 94350
rect 269738 94294 269808 94350
rect 269488 94226 269808 94294
rect 269488 94170 269558 94226
rect 269614 94170 269682 94226
rect 269738 94170 269808 94226
rect 269488 94102 269808 94170
rect 269488 94046 269558 94102
rect 269614 94046 269682 94102
rect 269738 94046 269808 94102
rect 269488 93978 269808 94046
rect 269488 93922 269558 93978
rect 269614 93922 269682 93978
rect 269738 93922 269808 93978
rect 269488 93888 269808 93922
rect 300208 94350 300528 94384
rect 300208 94294 300278 94350
rect 300334 94294 300402 94350
rect 300458 94294 300528 94350
rect 300208 94226 300528 94294
rect 300208 94170 300278 94226
rect 300334 94170 300402 94226
rect 300458 94170 300528 94226
rect 300208 94102 300528 94170
rect 300208 94046 300278 94102
rect 300334 94046 300402 94102
rect 300458 94046 300528 94102
rect 300208 93978 300528 94046
rect 300208 93922 300278 93978
rect 300334 93922 300402 93978
rect 300458 93922 300528 93978
rect 300208 93888 300528 93922
rect 330928 94350 331248 94384
rect 330928 94294 330998 94350
rect 331054 94294 331122 94350
rect 331178 94294 331248 94350
rect 330928 94226 331248 94294
rect 330928 94170 330998 94226
rect 331054 94170 331122 94226
rect 331178 94170 331248 94226
rect 330928 94102 331248 94170
rect 330928 94046 330998 94102
rect 331054 94046 331122 94102
rect 331178 94046 331248 94102
rect 330928 93978 331248 94046
rect 330928 93922 330998 93978
rect 331054 93922 331122 93978
rect 331178 93922 331248 93978
rect 330928 93888 331248 93922
rect 361648 94350 361968 94384
rect 361648 94294 361718 94350
rect 361774 94294 361842 94350
rect 361898 94294 361968 94350
rect 361648 94226 361968 94294
rect 361648 94170 361718 94226
rect 361774 94170 361842 94226
rect 361898 94170 361968 94226
rect 361648 94102 361968 94170
rect 361648 94046 361718 94102
rect 361774 94046 361842 94102
rect 361898 94046 361968 94102
rect 361648 93978 361968 94046
rect 361648 93922 361718 93978
rect 361774 93922 361842 93978
rect 361898 93922 361968 93978
rect 361648 93888 361968 93922
rect 392368 94350 392688 94384
rect 392368 94294 392438 94350
rect 392494 94294 392562 94350
rect 392618 94294 392688 94350
rect 392368 94226 392688 94294
rect 392368 94170 392438 94226
rect 392494 94170 392562 94226
rect 392618 94170 392688 94226
rect 392368 94102 392688 94170
rect 392368 94046 392438 94102
rect 392494 94046 392562 94102
rect 392618 94046 392688 94102
rect 392368 93978 392688 94046
rect 392368 93922 392438 93978
rect 392494 93922 392562 93978
rect 392618 93922 392688 93978
rect 392368 93888 392688 93922
rect 423088 94350 423408 94384
rect 423088 94294 423158 94350
rect 423214 94294 423282 94350
rect 423338 94294 423408 94350
rect 423088 94226 423408 94294
rect 423088 94170 423158 94226
rect 423214 94170 423282 94226
rect 423338 94170 423408 94226
rect 423088 94102 423408 94170
rect 423088 94046 423158 94102
rect 423214 94046 423282 94102
rect 423338 94046 423408 94102
rect 423088 93978 423408 94046
rect 423088 93922 423158 93978
rect 423214 93922 423282 93978
rect 423338 93922 423408 93978
rect 423088 93888 423408 93922
rect 453808 94350 454128 94384
rect 453808 94294 453878 94350
rect 453934 94294 454002 94350
rect 454058 94294 454128 94350
rect 453808 94226 454128 94294
rect 453808 94170 453878 94226
rect 453934 94170 454002 94226
rect 454058 94170 454128 94226
rect 453808 94102 454128 94170
rect 453808 94046 453878 94102
rect 453934 94046 454002 94102
rect 454058 94046 454128 94102
rect 453808 93978 454128 94046
rect 453808 93922 453878 93978
rect 453934 93922 454002 93978
rect 454058 93922 454128 93978
rect 453808 93888 454128 93922
rect 484528 94350 484848 94384
rect 484528 94294 484598 94350
rect 484654 94294 484722 94350
rect 484778 94294 484848 94350
rect 484528 94226 484848 94294
rect 484528 94170 484598 94226
rect 484654 94170 484722 94226
rect 484778 94170 484848 94226
rect 484528 94102 484848 94170
rect 484528 94046 484598 94102
rect 484654 94046 484722 94102
rect 484778 94046 484848 94102
rect 484528 93978 484848 94046
rect 484528 93922 484598 93978
rect 484654 93922 484722 93978
rect 484778 93922 484848 93978
rect 484528 93888 484848 93922
rect 515248 94350 515568 94384
rect 515248 94294 515318 94350
rect 515374 94294 515442 94350
rect 515498 94294 515568 94350
rect 515248 94226 515568 94294
rect 515248 94170 515318 94226
rect 515374 94170 515442 94226
rect 515498 94170 515568 94226
rect 515248 94102 515568 94170
rect 515248 94046 515318 94102
rect 515374 94046 515442 94102
rect 515498 94046 515568 94102
rect 515248 93978 515568 94046
rect 515248 93922 515318 93978
rect 515374 93922 515442 93978
rect 515498 93922 515568 93978
rect 515248 93888 515568 93922
rect 545968 94350 546288 94384
rect 545968 94294 546038 94350
rect 546094 94294 546162 94350
rect 546218 94294 546288 94350
rect 545968 94226 546288 94294
rect 545968 94170 546038 94226
rect 546094 94170 546162 94226
rect 546218 94170 546288 94226
rect 545968 94102 546288 94170
rect 545968 94046 546038 94102
rect 546094 94046 546162 94102
rect 546218 94046 546288 94102
rect 545968 93978 546288 94046
rect 545968 93922 546038 93978
rect 546094 93922 546162 93978
rect 546218 93922 546288 93978
rect 545968 93888 546288 93922
rect 561154 94350 561774 111922
rect 561154 94294 561250 94350
rect 561306 94294 561374 94350
rect 561430 94294 561498 94350
rect 561554 94294 561622 94350
rect 561678 94294 561774 94350
rect 561154 94226 561774 94294
rect 561154 94170 561250 94226
rect 561306 94170 561374 94226
rect 561430 94170 561498 94226
rect 561554 94170 561622 94226
rect 561678 94170 561774 94226
rect 561154 94102 561774 94170
rect 561154 94046 561250 94102
rect 561306 94046 561374 94102
rect 561430 94046 561498 94102
rect 561554 94046 561622 94102
rect 561678 94046 561774 94102
rect 561154 93978 561774 94046
rect 561154 93922 561250 93978
rect 561306 93922 561374 93978
rect 561430 93922 561498 93978
rect 561554 93922 561622 93978
rect 561678 93922 561774 93978
rect 131248 82350 131568 82384
rect 131248 82294 131318 82350
rect 131374 82294 131442 82350
rect 131498 82294 131568 82350
rect 131248 82226 131568 82294
rect 131248 82170 131318 82226
rect 131374 82170 131442 82226
rect 131498 82170 131568 82226
rect 131248 82102 131568 82170
rect 131248 82046 131318 82102
rect 131374 82046 131442 82102
rect 131498 82046 131568 82102
rect 131248 81978 131568 82046
rect 131248 81922 131318 81978
rect 131374 81922 131442 81978
rect 131498 81922 131568 81978
rect 131248 81888 131568 81922
rect 161968 82350 162288 82384
rect 161968 82294 162038 82350
rect 162094 82294 162162 82350
rect 162218 82294 162288 82350
rect 161968 82226 162288 82294
rect 161968 82170 162038 82226
rect 162094 82170 162162 82226
rect 162218 82170 162288 82226
rect 161968 82102 162288 82170
rect 161968 82046 162038 82102
rect 162094 82046 162162 82102
rect 162218 82046 162288 82102
rect 161968 81978 162288 82046
rect 161968 81922 162038 81978
rect 162094 81922 162162 81978
rect 162218 81922 162288 81978
rect 161968 81888 162288 81922
rect 192688 82350 193008 82384
rect 192688 82294 192758 82350
rect 192814 82294 192882 82350
rect 192938 82294 193008 82350
rect 192688 82226 193008 82294
rect 192688 82170 192758 82226
rect 192814 82170 192882 82226
rect 192938 82170 193008 82226
rect 192688 82102 193008 82170
rect 192688 82046 192758 82102
rect 192814 82046 192882 82102
rect 192938 82046 193008 82102
rect 192688 81978 193008 82046
rect 192688 81922 192758 81978
rect 192814 81922 192882 81978
rect 192938 81922 193008 81978
rect 192688 81888 193008 81922
rect 223408 82350 223728 82384
rect 223408 82294 223478 82350
rect 223534 82294 223602 82350
rect 223658 82294 223728 82350
rect 223408 82226 223728 82294
rect 223408 82170 223478 82226
rect 223534 82170 223602 82226
rect 223658 82170 223728 82226
rect 223408 82102 223728 82170
rect 223408 82046 223478 82102
rect 223534 82046 223602 82102
rect 223658 82046 223728 82102
rect 223408 81978 223728 82046
rect 223408 81922 223478 81978
rect 223534 81922 223602 81978
rect 223658 81922 223728 81978
rect 223408 81888 223728 81922
rect 254128 82350 254448 82384
rect 254128 82294 254198 82350
rect 254254 82294 254322 82350
rect 254378 82294 254448 82350
rect 254128 82226 254448 82294
rect 254128 82170 254198 82226
rect 254254 82170 254322 82226
rect 254378 82170 254448 82226
rect 254128 82102 254448 82170
rect 254128 82046 254198 82102
rect 254254 82046 254322 82102
rect 254378 82046 254448 82102
rect 254128 81978 254448 82046
rect 254128 81922 254198 81978
rect 254254 81922 254322 81978
rect 254378 81922 254448 81978
rect 254128 81888 254448 81922
rect 284848 82350 285168 82384
rect 284848 82294 284918 82350
rect 284974 82294 285042 82350
rect 285098 82294 285168 82350
rect 284848 82226 285168 82294
rect 284848 82170 284918 82226
rect 284974 82170 285042 82226
rect 285098 82170 285168 82226
rect 284848 82102 285168 82170
rect 284848 82046 284918 82102
rect 284974 82046 285042 82102
rect 285098 82046 285168 82102
rect 284848 81978 285168 82046
rect 284848 81922 284918 81978
rect 284974 81922 285042 81978
rect 285098 81922 285168 81978
rect 284848 81888 285168 81922
rect 315568 82350 315888 82384
rect 315568 82294 315638 82350
rect 315694 82294 315762 82350
rect 315818 82294 315888 82350
rect 315568 82226 315888 82294
rect 315568 82170 315638 82226
rect 315694 82170 315762 82226
rect 315818 82170 315888 82226
rect 315568 82102 315888 82170
rect 315568 82046 315638 82102
rect 315694 82046 315762 82102
rect 315818 82046 315888 82102
rect 315568 81978 315888 82046
rect 315568 81922 315638 81978
rect 315694 81922 315762 81978
rect 315818 81922 315888 81978
rect 315568 81888 315888 81922
rect 346288 82350 346608 82384
rect 346288 82294 346358 82350
rect 346414 82294 346482 82350
rect 346538 82294 346608 82350
rect 346288 82226 346608 82294
rect 346288 82170 346358 82226
rect 346414 82170 346482 82226
rect 346538 82170 346608 82226
rect 346288 82102 346608 82170
rect 346288 82046 346358 82102
rect 346414 82046 346482 82102
rect 346538 82046 346608 82102
rect 346288 81978 346608 82046
rect 346288 81922 346358 81978
rect 346414 81922 346482 81978
rect 346538 81922 346608 81978
rect 346288 81888 346608 81922
rect 377008 82350 377328 82384
rect 377008 82294 377078 82350
rect 377134 82294 377202 82350
rect 377258 82294 377328 82350
rect 377008 82226 377328 82294
rect 377008 82170 377078 82226
rect 377134 82170 377202 82226
rect 377258 82170 377328 82226
rect 377008 82102 377328 82170
rect 377008 82046 377078 82102
rect 377134 82046 377202 82102
rect 377258 82046 377328 82102
rect 377008 81978 377328 82046
rect 377008 81922 377078 81978
rect 377134 81922 377202 81978
rect 377258 81922 377328 81978
rect 377008 81888 377328 81922
rect 407728 82350 408048 82384
rect 407728 82294 407798 82350
rect 407854 82294 407922 82350
rect 407978 82294 408048 82350
rect 407728 82226 408048 82294
rect 407728 82170 407798 82226
rect 407854 82170 407922 82226
rect 407978 82170 408048 82226
rect 407728 82102 408048 82170
rect 407728 82046 407798 82102
rect 407854 82046 407922 82102
rect 407978 82046 408048 82102
rect 407728 81978 408048 82046
rect 407728 81922 407798 81978
rect 407854 81922 407922 81978
rect 407978 81922 408048 81978
rect 407728 81888 408048 81922
rect 438448 82350 438768 82384
rect 438448 82294 438518 82350
rect 438574 82294 438642 82350
rect 438698 82294 438768 82350
rect 438448 82226 438768 82294
rect 438448 82170 438518 82226
rect 438574 82170 438642 82226
rect 438698 82170 438768 82226
rect 438448 82102 438768 82170
rect 438448 82046 438518 82102
rect 438574 82046 438642 82102
rect 438698 82046 438768 82102
rect 438448 81978 438768 82046
rect 438448 81922 438518 81978
rect 438574 81922 438642 81978
rect 438698 81922 438768 81978
rect 438448 81888 438768 81922
rect 469168 82350 469488 82384
rect 469168 82294 469238 82350
rect 469294 82294 469362 82350
rect 469418 82294 469488 82350
rect 469168 82226 469488 82294
rect 469168 82170 469238 82226
rect 469294 82170 469362 82226
rect 469418 82170 469488 82226
rect 469168 82102 469488 82170
rect 469168 82046 469238 82102
rect 469294 82046 469362 82102
rect 469418 82046 469488 82102
rect 469168 81978 469488 82046
rect 469168 81922 469238 81978
rect 469294 81922 469362 81978
rect 469418 81922 469488 81978
rect 469168 81888 469488 81922
rect 499888 82350 500208 82384
rect 499888 82294 499958 82350
rect 500014 82294 500082 82350
rect 500138 82294 500208 82350
rect 499888 82226 500208 82294
rect 499888 82170 499958 82226
rect 500014 82170 500082 82226
rect 500138 82170 500208 82226
rect 499888 82102 500208 82170
rect 499888 82046 499958 82102
rect 500014 82046 500082 82102
rect 500138 82046 500208 82102
rect 499888 81978 500208 82046
rect 499888 81922 499958 81978
rect 500014 81922 500082 81978
rect 500138 81922 500208 81978
rect 499888 81888 500208 81922
rect 530608 82350 530928 82384
rect 530608 82294 530678 82350
rect 530734 82294 530802 82350
rect 530858 82294 530928 82350
rect 530608 82226 530928 82294
rect 530608 82170 530678 82226
rect 530734 82170 530802 82226
rect 530858 82170 530928 82226
rect 530608 82102 530928 82170
rect 530608 82046 530678 82102
rect 530734 82046 530802 82102
rect 530858 82046 530928 82102
rect 530608 81978 530928 82046
rect 530608 81922 530678 81978
rect 530734 81922 530802 81978
rect 530858 81922 530928 81978
rect 530608 81888 530928 81922
rect 111154 76294 111250 76350
rect 111306 76294 111374 76350
rect 111430 76294 111498 76350
rect 111554 76294 111622 76350
rect 111678 76294 111774 76350
rect 111154 76226 111774 76294
rect 111154 76170 111250 76226
rect 111306 76170 111374 76226
rect 111430 76170 111498 76226
rect 111554 76170 111622 76226
rect 111678 76170 111774 76226
rect 111154 76102 111774 76170
rect 111154 76046 111250 76102
rect 111306 76046 111374 76102
rect 111430 76046 111498 76102
rect 111554 76046 111622 76102
rect 111678 76046 111774 76102
rect 111154 75978 111774 76046
rect 111154 75922 111250 75978
rect 111306 75922 111374 75978
rect 111430 75922 111498 75978
rect 111554 75922 111622 75978
rect 111678 75922 111774 75978
rect 96874 64294 96970 64350
rect 97026 64294 97094 64350
rect 97150 64294 97218 64350
rect 97274 64294 97342 64350
rect 97398 64294 97494 64350
rect 96874 64226 97494 64294
rect 96874 64170 96970 64226
rect 97026 64170 97094 64226
rect 97150 64170 97218 64226
rect 97274 64170 97342 64226
rect 97398 64170 97494 64226
rect 96874 64102 97494 64170
rect 96874 64046 96970 64102
rect 97026 64046 97094 64102
rect 97150 64046 97218 64102
rect 97274 64046 97342 64102
rect 97398 64046 97494 64102
rect 96874 63978 97494 64046
rect 96874 63922 96970 63978
rect 97026 63922 97094 63978
rect 97150 63922 97218 63978
rect 97274 63922 97342 63978
rect 97398 63922 97494 63978
rect 96874 46350 97494 63922
rect 100528 64350 100848 64384
rect 100528 64294 100598 64350
rect 100654 64294 100722 64350
rect 100778 64294 100848 64350
rect 100528 64226 100848 64294
rect 100528 64170 100598 64226
rect 100654 64170 100722 64226
rect 100778 64170 100848 64226
rect 100528 64102 100848 64170
rect 100528 64046 100598 64102
rect 100654 64046 100722 64102
rect 100778 64046 100848 64102
rect 100528 63978 100848 64046
rect 100528 63922 100598 63978
rect 100654 63922 100722 63978
rect 100778 63922 100848 63978
rect 100528 63888 100848 63922
rect 111154 58350 111774 75922
rect 115888 76350 116208 76384
rect 115888 76294 115958 76350
rect 116014 76294 116082 76350
rect 116138 76294 116208 76350
rect 115888 76226 116208 76294
rect 115888 76170 115958 76226
rect 116014 76170 116082 76226
rect 116138 76170 116208 76226
rect 115888 76102 116208 76170
rect 115888 76046 115958 76102
rect 116014 76046 116082 76102
rect 116138 76046 116208 76102
rect 115888 75978 116208 76046
rect 115888 75922 115958 75978
rect 116014 75922 116082 75978
rect 116138 75922 116208 75978
rect 115888 75888 116208 75922
rect 146608 76350 146928 76384
rect 146608 76294 146678 76350
rect 146734 76294 146802 76350
rect 146858 76294 146928 76350
rect 146608 76226 146928 76294
rect 146608 76170 146678 76226
rect 146734 76170 146802 76226
rect 146858 76170 146928 76226
rect 146608 76102 146928 76170
rect 146608 76046 146678 76102
rect 146734 76046 146802 76102
rect 146858 76046 146928 76102
rect 146608 75978 146928 76046
rect 146608 75922 146678 75978
rect 146734 75922 146802 75978
rect 146858 75922 146928 75978
rect 146608 75888 146928 75922
rect 177328 76350 177648 76384
rect 177328 76294 177398 76350
rect 177454 76294 177522 76350
rect 177578 76294 177648 76350
rect 177328 76226 177648 76294
rect 177328 76170 177398 76226
rect 177454 76170 177522 76226
rect 177578 76170 177648 76226
rect 177328 76102 177648 76170
rect 177328 76046 177398 76102
rect 177454 76046 177522 76102
rect 177578 76046 177648 76102
rect 177328 75978 177648 76046
rect 177328 75922 177398 75978
rect 177454 75922 177522 75978
rect 177578 75922 177648 75978
rect 177328 75888 177648 75922
rect 208048 76350 208368 76384
rect 208048 76294 208118 76350
rect 208174 76294 208242 76350
rect 208298 76294 208368 76350
rect 208048 76226 208368 76294
rect 208048 76170 208118 76226
rect 208174 76170 208242 76226
rect 208298 76170 208368 76226
rect 208048 76102 208368 76170
rect 208048 76046 208118 76102
rect 208174 76046 208242 76102
rect 208298 76046 208368 76102
rect 208048 75978 208368 76046
rect 208048 75922 208118 75978
rect 208174 75922 208242 75978
rect 208298 75922 208368 75978
rect 208048 75888 208368 75922
rect 238768 76350 239088 76384
rect 238768 76294 238838 76350
rect 238894 76294 238962 76350
rect 239018 76294 239088 76350
rect 238768 76226 239088 76294
rect 238768 76170 238838 76226
rect 238894 76170 238962 76226
rect 239018 76170 239088 76226
rect 238768 76102 239088 76170
rect 238768 76046 238838 76102
rect 238894 76046 238962 76102
rect 239018 76046 239088 76102
rect 238768 75978 239088 76046
rect 238768 75922 238838 75978
rect 238894 75922 238962 75978
rect 239018 75922 239088 75978
rect 238768 75888 239088 75922
rect 269488 76350 269808 76384
rect 269488 76294 269558 76350
rect 269614 76294 269682 76350
rect 269738 76294 269808 76350
rect 269488 76226 269808 76294
rect 269488 76170 269558 76226
rect 269614 76170 269682 76226
rect 269738 76170 269808 76226
rect 269488 76102 269808 76170
rect 269488 76046 269558 76102
rect 269614 76046 269682 76102
rect 269738 76046 269808 76102
rect 269488 75978 269808 76046
rect 269488 75922 269558 75978
rect 269614 75922 269682 75978
rect 269738 75922 269808 75978
rect 269488 75888 269808 75922
rect 300208 76350 300528 76384
rect 300208 76294 300278 76350
rect 300334 76294 300402 76350
rect 300458 76294 300528 76350
rect 300208 76226 300528 76294
rect 300208 76170 300278 76226
rect 300334 76170 300402 76226
rect 300458 76170 300528 76226
rect 300208 76102 300528 76170
rect 300208 76046 300278 76102
rect 300334 76046 300402 76102
rect 300458 76046 300528 76102
rect 300208 75978 300528 76046
rect 300208 75922 300278 75978
rect 300334 75922 300402 75978
rect 300458 75922 300528 75978
rect 300208 75888 300528 75922
rect 330928 76350 331248 76384
rect 330928 76294 330998 76350
rect 331054 76294 331122 76350
rect 331178 76294 331248 76350
rect 330928 76226 331248 76294
rect 330928 76170 330998 76226
rect 331054 76170 331122 76226
rect 331178 76170 331248 76226
rect 330928 76102 331248 76170
rect 330928 76046 330998 76102
rect 331054 76046 331122 76102
rect 331178 76046 331248 76102
rect 330928 75978 331248 76046
rect 330928 75922 330998 75978
rect 331054 75922 331122 75978
rect 331178 75922 331248 75978
rect 330928 75888 331248 75922
rect 361648 76350 361968 76384
rect 361648 76294 361718 76350
rect 361774 76294 361842 76350
rect 361898 76294 361968 76350
rect 361648 76226 361968 76294
rect 361648 76170 361718 76226
rect 361774 76170 361842 76226
rect 361898 76170 361968 76226
rect 361648 76102 361968 76170
rect 361648 76046 361718 76102
rect 361774 76046 361842 76102
rect 361898 76046 361968 76102
rect 361648 75978 361968 76046
rect 361648 75922 361718 75978
rect 361774 75922 361842 75978
rect 361898 75922 361968 75978
rect 361648 75888 361968 75922
rect 392368 76350 392688 76384
rect 392368 76294 392438 76350
rect 392494 76294 392562 76350
rect 392618 76294 392688 76350
rect 392368 76226 392688 76294
rect 392368 76170 392438 76226
rect 392494 76170 392562 76226
rect 392618 76170 392688 76226
rect 392368 76102 392688 76170
rect 392368 76046 392438 76102
rect 392494 76046 392562 76102
rect 392618 76046 392688 76102
rect 392368 75978 392688 76046
rect 392368 75922 392438 75978
rect 392494 75922 392562 75978
rect 392618 75922 392688 75978
rect 392368 75888 392688 75922
rect 423088 76350 423408 76384
rect 423088 76294 423158 76350
rect 423214 76294 423282 76350
rect 423338 76294 423408 76350
rect 423088 76226 423408 76294
rect 423088 76170 423158 76226
rect 423214 76170 423282 76226
rect 423338 76170 423408 76226
rect 423088 76102 423408 76170
rect 423088 76046 423158 76102
rect 423214 76046 423282 76102
rect 423338 76046 423408 76102
rect 423088 75978 423408 76046
rect 423088 75922 423158 75978
rect 423214 75922 423282 75978
rect 423338 75922 423408 75978
rect 423088 75888 423408 75922
rect 453808 76350 454128 76384
rect 453808 76294 453878 76350
rect 453934 76294 454002 76350
rect 454058 76294 454128 76350
rect 453808 76226 454128 76294
rect 453808 76170 453878 76226
rect 453934 76170 454002 76226
rect 454058 76170 454128 76226
rect 453808 76102 454128 76170
rect 453808 76046 453878 76102
rect 453934 76046 454002 76102
rect 454058 76046 454128 76102
rect 453808 75978 454128 76046
rect 453808 75922 453878 75978
rect 453934 75922 454002 75978
rect 454058 75922 454128 75978
rect 453808 75888 454128 75922
rect 484528 76350 484848 76384
rect 484528 76294 484598 76350
rect 484654 76294 484722 76350
rect 484778 76294 484848 76350
rect 484528 76226 484848 76294
rect 484528 76170 484598 76226
rect 484654 76170 484722 76226
rect 484778 76170 484848 76226
rect 484528 76102 484848 76170
rect 484528 76046 484598 76102
rect 484654 76046 484722 76102
rect 484778 76046 484848 76102
rect 484528 75978 484848 76046
rect 484528 75922 484598 75978
rect 484654 75922 484722 75978
rect 484778 75922 484848 75978
rect 484528 75888 484848 75922
rect 515248 76350 515568 76384
rect 515248 76294 515318 76350
rect 515374 76294 515442 76350
rect 515498 76294 515568 76350
rect 515248 76226 515568 76294
rect 515248 76170 515318 76226
rect 515374 76170 515442 76226
rect 515498 76170 515568 76226
rect 515248 76102 515568 76170
rect 515248 76046 515318 76102
rect 515374 76046 515442 76102
rect 515498 76046 515568 76102
rect 515248 75978 515568 76046
rect 515248 75922 515318 75978
rect 515374 75922 515442 75978
rect 515498 75922 515568 75978
rect 515248 75888 515568 75922
rect 545968 76350 546288 76384
rect 545968 76294 546038 76350
rect 546094 76294 546162 76350
rect 546218 76294 546288 76350
rect 545968 76226 546288 76294
rect 545968 76170 546038 76226
rect 546094 76170 546162 76226
rect 546218 76170 546288 76226
rect 545968 76102 546288 76170
rect 545968 76046 546038 76102
rect 546094 76046 546162 76102
rect 546218 76046 546288 76102
rect 545968 75978 546288 76046
rect 545968 75922 546038 75978
rect 546094 75922 546162 75978
rect 546218 75922 546288 75978
rect 545968 75888 546288 75922
rect 561154 76350 561774 93922
rect 561154 76294 561250 76350
rect 561306 76294 561374 76350
rect 561430 76294 561498 76350
rect 561554 76294 561622 76350
rect 561678 76294 561774 76350
rect 561154 76226 561774 76294
rect 561154 76170 561250 76226
rect 561306 76170 561374 76226
rect 561430 76170 561498 76226
rect 561554 76170 561622 76226
rect 561678 76170 561774 76226
rect 561154 76102 561774 76170
rect 561154 76046 561250 76102
rect 561306 76046 561374 76102
rect 561430 76046 561498 76102
rect 561554 76046 561622 76102
rect 561678 76046 561774 76102
rect 561154 75978 561774 76046
rect 561154 75922 561250 75978
rect 561306 75922 561374 75978
rect 561430 75922 561498 75978
rect 561554 75922 561622 75978
rect 561678 75922 561774 75978
rect 131248 64350 131568 64384
rect 131248 64294 131318 64350
rect 131374 64294 131442 64350
rect 131498 64294 131568 64350
rect 131248 64226 131568 64294
rect 131248 64170 131318 64226
rect 131374 64170 131442 64226
rect 131498 64170 131568 64226
rect 131248 64102 131568 64170
rect 131248 64046 131318 64102
rect 131374 64046 131442 64102
rect 131498 64046 131568 64102
rect 131248 63978 131568 64046
rect 131248 63922 131318 63978
rect 131374 63922 131442 63978
rect 131498 63922 131568 63978
rect 131248 63888 131568 63922
rect 161968 64350 162288 64384
rect 161968 64294 162038 64350
rect 162094 64294 162162 64350
rect 162218 64294 162288 64350
rect 161968 64226 162288 64294
rect 161968 64170 162038 64226
rect 162094 64170 162162 64226
rect 162218 64170 162288 64226
rect 161968 64102 162288 64170
rect 161968 64046 162038 64102
rect 162094 64046 162162 64102
rect 162218 64046 162288 64102
rect 161968 63978 162288 64046
rect 161968 63922 162038 63978
rect 162094 63922 162162 63978
rect 162218 63922 162288 63978
rect 161968 63888 162288 63922
rect 192688 64350 193008 64384
rect 192688 64294 192758 64350
rect 192814 64294 192882 64350
rect 192938 64294 193008 64350
rect 192688 64226 193008 64294
rect 192688 64170 192758 64226
rect 192814 64170 192882 64226
rect 192938 64170 193008 64226
rect 192688 64102 193008 64170
rect 192688 64046 192758 64102
rect 192814 64046 192882 64102
rect 192938 64046 193008 64102
rect 192688 63978 193008 64046
rect 192688 63922 192758 63978
rect 192814 63922 192882 63978
rect 192938 63922 193008 63978
rect 192688 63888 193008 63922
rect 223408 64350 223728 64384
rect 223408 64294 223478 64350
rect 223534 64294 223602 64350
rect 223658 64294 223728 64350
rect 223408 64226 223728 64294
rect 223408 64170 223478 64226
rect 223534 64170 223602 64226
rect 223658 64170 223728 64226
rect 223408 64102 223728 64170
rect 223408 64046 223478 64102
rect 223534 64046 223602 64102
rect 223658 64046 223728 64102
rect 223408 63978 223728 64046
rect 223408 63922 223478 63978
rect 223534 63922 223602 63978
rect 223658 63922 223728 63978
rect 223408 63888 223728 63922
rect 254128 64350 254448 64384
rect 254128 64294 254198 64350
rect 254254 64294 254322 64350
rect 254378 64294 254448 64350
rect 254128 64226 254448 64294
rect 254128 64170 254198 64226
rect 254254 64170 254322 64226
rect 254378 64170 254448 64226
rect 254128 64102 254448 64170
rect 254128 64046 254198 64102
rect 254254 64046 254322 64102
rect 254378 64046 254448 64102
rect 254128 63978 254448 64046
rect 254128 63922 254198 63978
rect 254254 63922 254322 63978
rect 254378 63922 254448 63978
rect 254128 63888 254448 63922
rect 284848 64350 285168 64384
rect 284848 64294 284918 64350
rect 284974 64294 285042 64350
rect 285098 64294 285168 64350
rect 284848 64226 285168 64294
rect 284848 64170 284918 64226
rect 284974 64170 285042 64226
rect 285098 64170 285168 64226
rect 284848 64102 285168 64170
rect 284848 64046 284918 64102
rect 284974 64046 285042 64102
rect 285098 64046 285168 64102
rect 284848 63978 285168 64046
rect 284848 63922 284918 63978
rect 284974 63922 285042 63978
rect 285098 63922 285168 63978
rect 284848 63888 285168 63922
rect 315568 64350 315888 64384
rect 315568 64294 315638 64350
rect 315694 64294 315762 64350
rect 315818 64294 315888 64350
rect 315568 64226 315888 64294
rect 315568 64170 315638 64226
rect 315694 64170 315762 64226
rect 315818 64170 315888 64226
rect 315568 64102 315888 64170
rect 315568 64046 315638 64102
rect 315694 64046 315762 64102
rect 315818 64046 315888 64102
rect 315568 63978 315888 64046
rect 315568 63922 315638 63978
rect 315694 63922 315762 63978
rect 315818 63922 315888 63978
rect 315568 63888 315888 63922
rect 346288 64350 346608 64384
rect 346288 64294 346358 64350
rect 346414 64294 346482 64350
rect 346538 64294 346608 64350
rect 346288 64226 346608 64294
rect 346288 64170 346358 64226
rect 346414 64170 346482 64226
rect 346538 64170 346608 64226
rect 346288 64102 346608 64170
rect 346288 64046 346358 64102
rect 346414 64046 346482 64102
rect 346538 64046 346608 64102
rect 346288 63978 346608 64046
rect 346288 63922 346358 63978
rect 346414 63922 346482 63978
rect 346538 63922 346608 63978
rect 346288 63888 346608 63922
rect 377008 64350 377328 64384
rect 377008 64294 377078 64350
rect 377134 64294 377202 64350
rect 377258 64294 377328 64350
rect 377008 64226 377328 64294
rect 377008 64170 377078 64226
rect 377134 64170 377202 64226
rect 377258 64170 377328 64226
rect 377008 64102 377328 64170
rect 377008 64046 377078 64102
rect 377134 64046 377202 64102
rect 377258 64046 377328 64102
rect 377008 63978 377328 64046
rect 377008 63922 377078 63978
rect 377134 63922 377202 63978
rect 377258 63922 377328 63978
rect 377008 63888 377328 63922
rect 407728 64350 408048 64384
rect 407728 64294 407798 64350
rect 407854 64294 407922 64350
rect 407978 64294 408048 64350
rect 407728 64226 408048 64294
rect 407728 64170 407798 64226
rect 407854 64170 407922 64226
rect 407978 64170 408048 64226
rect 407728 64102 408048 64170
rect 407728 64046 407798 64102
rect 407854 64046 407922 64102
rect 407978 64046 408048 64102
rect 407728 63978 408048 64046
rect 407728 63922 407798 63978
rect 407854 63922 407922 63978
rect 407978 63922 408048 63978
rect 407728 63888 408048 63922
rect 438448 64350 438768 64384
rect 438448 64294 438518 64350
rect 438574 64294 438642 64350
rect 438698 64294 438768 64350
rect 438448 64226 438768 64294
rect 438448 64170 438518 64226
rect 438574 64170 438642 64226
rect 438698 64170 438768 64226
rect 438448 64102 438768 64170
rect 438448 64046 438518 64102
rect 438574 64046 438642 64102
rect 438698 64046 438768 64102
rect 438448 63978 438768 64046
rect 438448 63922 438518 63978
rect 438574 63922 438642 63978
rect 438698 63922 438768 63978
rect 438448 63888 438768 63922
rect 469168 64350 469488 64384
rect 469168 64294 469238 64350
rect 469294 64294 469362 64350
rect 469418 64294 469488 64350
rect 469168 64226 469488 64294
rect 469168 64170 469238 64226
rect 469294 64170 469362 64226
rect 469418 64170 469488 64226
rect 469168 64102 469488 64170
rect 469168 64046 469238 64102
rect 469294 64046 469362 64102
rect 469418 64046 469488 64102
rect 469168 63978 469488 64046
rect 469168 63922 469238 63978
rect 469294 63922 469362 63978
rect 469418 63922 469488 63978
rect 469168 63888 469488 63922
rect 499888 64350 500208 64384
rect 499888 64294 499958 64350
rect 500014 64294 500082 64350
rect 500138 64294 500208 64350
rect 499888 64226 500208 64294
rect 499888 64170 499958 64226
rect 500014 64170 500082 64226
rect 500138 64170 500208 64226
rect 499888 64102 500208 64170
rect 499888 64046 499958 64102
rect 500014 64046 500082 64102
rect 500138 64046 500208 64102
rect 499888 63978 500208 64046
rect 499888 63922 499958 63978
rect 500014 63922 500082 63978
rect 500138 63922 500208 63978
rect 499888 63888 500208 63922
rect 530608 64350 530928 64384
rect 530608 64294 530678 64350
rect 530734 64294 530802 64350
rect 530858 64294 530928 64350
rect 530608 64226 530928 64294
rect 530608 64170 530678 64226
rect 530734 64170 530802 64226
rect 530858 64170 530928 64226
rect 530608 64102 530928 64170
rect 530608 64046 530678 64102
rect 530734 64046 530802 64102
rect 530858 64046 530928 64102
rect 530608 63978 530928 64046
rect 530608 63922 530678 63978
rect 530734 63922 530802 63978
rect 530858 63922 530928 63978
rect 530608 63888 530928 63922
rect 111154 58294 111250 58350
rect 111306 58294 111374 58350
rect 111430 58294 111498 58350
rect 111554 58294 111622 58350
rect 111678 58294 111774 58350
rect 111154 58226 111774 58294
rect 111154 58170 111250 58226
rect 111306 58170 111374 58226
rect 111430 58170 111498 58226
rect 111554 58170 111622 58226
rect 111678 58170 111774 58226
rect 111154 58102 111774 58170
rect 111154 58046 111250 58102
rect 111306 58046 111374 58102
rect 111430 58046 111498 58102
rect 111554 58046 111622 58102
rect 111678 58046 111774 58102
rect 111154 57978 111774 58046
rect 111154 57922 111250 57978
rect 111306 57922 111374 57978
rect 111430 57922 111498 57978
rect 111554 57922 111622 57978
rect 111678 57922 111774 57978
rect 96874 46294 96970 46350
rect 97026 46294 97094 46350
rect 97150 46294 97218 46350
rect 97274 46294 97342 46350
rect 97398 46294 97494 46350
rect 96874 46226 97494 46294
rect 96874 46170 96970 46226
rect 97026 46170 97094 46226
rect 97150 46170 97218 46226
rect 97274 46170 97342 46226
rect 97398 46170 97494 46226
rect 96874 46102 97494 46170
rect 96874 46046 96970 46102
rect 97026 46046 97094 46102
rect 97150 46046 97218 46102
rect 97274 46046 97342 46102
rect 97398 46046 97494 46102
rect 96874 45978 97494 46046
rect 96874 45922 96970 45978
rect 97026 45922 97094 45978
rect 97150 45922 97218 45978
rect 97274 45922 97342 45978
rect 97398 45922 97494 45978
rect 96874 28350 97494 45922
rect 100528 46350 100848 46384
rect 100528 46294 100598 46350
rect 100654 46294 100722 46350
rect 100778 46294 100848 46350
rect 100528 46226 100848 46294
rect 100528 46170 100598 46226
rect 100654 46170 100722 46226
rect 100778 46170 100848 46226
rect 100528 46102 100848 46170
rect 100528 46046 100598 46102
rect 100654 46046 100722 46102
rect 100778 46046 100848 46102
rect 100528 45978 100848 46046
rect 100528 45922 100598 45978
rect 100654 45922 100722 45978
rect 100778 45922 100848 45978
rect 100528 45888 100848 45922
rect 96874 28294 96970 28350
rect 97026 28294 97094 28350
rect 97150 28294 97218 28350
rect 97274 28294 97342 28350
rect 97398 28294 97494 28350
rect 96874 28226 97494 28294
rect 96874 28170 96970 28226
rect 97026 28170 97094 28226
rect 97150 28170 97218 28226
rect 97274 28170 97342 28226
rect 97398 28170 97494 28226
rect 96874 28102 97494 28170
rect 96874 28046 96970 28102
rect 97026 28046 97094 28102
rect 97150 28046 97218 28102
rect 97274 28046 97342 28102
rect 97398 28046 97494 28102
rect 96874 27978 97494 28046
rect 96874 27922 96970 27978
rect 97026 27922 97094 27978
rect 97150 27922 97218 27978
rect 97274 27922 97342 27978
rect 97398 27922 97494 27978
rect 96874 10350 97494 27922
rect 96874 10294 96970 10350
rect 97026 10294 97094 10350
rect 97150 10294 97218 10350
rect 97274 10294 97342 10350
rect 97398 10294 97494 10350
rect 96874 10226 97494 10294
rect 96874 10170 96970 10226
rect 97026 10170 97094 10226
rect 97150 10170 97218 10226
rect 97274 10170 97342 10226
rect 97398 10170 97494 10226
rect 96874 10102 97494 10170
rect 96874 10046 96970 10102
rect 97026 10046 97094 10102
rect 97150 10046 97218 10102
rect 97274 10046 97342 10102
rect 97398 10046 97494 10102
rect 96874 9978 97494 10046
rect 96874 9922 96970 9978
rect 97026 9922 97094 9978
rect 97150 9922 97218 9978
rect 97274 9922 97342 9978
rect 97398 9922 97494 9978
rect 96874 -1120 97494 9922
rect 96874 -1176 96970 -1120
rect 97026 -1176 97094 -1120
rect 97150 -1176 97218 -1120
rect 97274 -1176 97342 -1120
rect 97398 -1176 97494 -1120
rect 96874 -1244 97494 -1176
rect 96874 -1300 96970 -1244
rect 97026 -1300 97094 -1244
rect 97150 -1300 97218 -1244
rect 97274 -1300 97342 -1244
rect 97398 -1300 97494 -1244
rect 96874 -1368 97494 -1300
rect 96874 -1424 96970 -1368
rect 97026 -1424 97094 -1368
rect 97150 -1424 97218 -1368
rect 97274 -1424 97342 -1368
rect 97398 -1424 97494 -1368
rect 96874 -1492 97494 -1424
rect 96874 -1548 96970 -1492
rect 97026 -1548 97094 -1492
rect 97150 -1548 97218 -1492
rect 97274 -1548 97342 -1492
rect 97398 -1548 97494 -1492
rect 96874 -1644 97494 -1548
rect 111154 40350 111774 57922
rect 115888 58350 116208 58384
rect 115888 58294 115958 58350
rect 116014 58294 116082 58350
rect 116138 58294 116208 58350
rect 115888 58226 116208 58294
rect 115888 58170 115958 58226
rect 116014 58170 116082 58226
rect 116138 58170 116208 58226
rect 115888 58102 116208 58170
rect 115888 58046 115958 58102
rect 116014 58046 116082 58102
rect 116138 58046 116208 58102
rect 115888 57978 116208 58046
rect 115888 57922 115958 57978
rect 116014 57922 116082 57978
rect 116138 57922 116208 57978
rect 115888 57888 116208 57922
rect 146608 58350 146928 58384
rect 146608 58294 146678 58350
rect 146734 58294 146802 58350
rect 146858 58294 146928 58350
rect 146608 58226 146928 58294
rect 146608 58170 146678 58226
rect 146734 58170 146802 58226
rect 146858 58170 146928 58226
rect 146608 58102 146928 58170
rect 146608 58046 146678 58102
rect 146734 58046 146802 58102
rect 146858 58046 146928 58102
rect 146608 57978 146928 58046
rect 146608 57922 146678 57978
rect 146734 57922 146802 57978
rect 146858 57922 146928 57978
rect 146608 57888 146928 57922
rect 177328 58350 177648 58384
rect 177328 58294 177398 58350
rect 177454 58294 177522 58350
rect 177578 58294 177648 58350
rect 177328 58226 177648 58294
rect 177328 58170 177398 58226
rect 177454 58170 177522 58226
rect 177578 58170 177648 58226
rect 177328 58102 177648 58170
rect 177328 58046 177398 58102
rect 177454 58046 177522 58102
rect 177578 58046 177648 58102
rect 177328 57978 177648 58046
rect 177328 57922 177398 57978
rect 177454 57922 177522 57978
rect 177578 57922 177648 57978
rect 177328 57888 177648 57922
rect 208048 58350 208368 58384
rect 208048 58294 208118 58350
rect 208174 58294 208242 58350
rect 208298 58294 208368 58350
rect 208048 58226 208368 58294
rect 208048 58170 208118 58226
rect 208174 58170 208242 58226
rect 208298 58170 208368 58226
rect 208048 58102 208368 58170
rect 208048 58046 208118 58102
rect 208174 58046 208242 58102
rect 208298 58046 208368 58102
rect 208048 57978 208368 58046
rect 208048 57922 208118 57978
rect 208174 57922 208242 57978
rect 208298 57922 208368 57978
rect 208048 57888 208368 57922
rect 238768 58350 239088 58384
rect 238768 58294 238838 58350
rect 238894 58294 238962 58350
rect 239018 58294 239088 58350
rect 238768 58226 239088 58294
rect 238768 58170 238838 58226
rect 238894 58170 238962 58226
rect 239018 58170 239088 58226
rect 238768 58102 239088 58170
rect 238768 58046 238838 58102
rect 238894 58046 238962 58102
rect 239018 58046 239088 58102
rect 238768 57978 239088 58046
rect 238768 57922 238838 57978
rect 238894 57922 238962 57978
rect 239018 57922 239088 57978
rect 238768 57888 239088 57922
rect 269488 58350 269808 58384
rect 269488 58294 269558 58350
rect 269614 58294 269682 58350
rect 269738 58294 269808 58350
rect 269488 58226 269808 58294
rect 269488 58170 269558 58226
rect 269614 58170 269682 58226
rect 269738 58170 269808 58226
rect 269488 58102 269808 58170
rect 269488 58046 269558 58102
rect 269614 58046 269682 58102
rect 269738 58046 269808 58102
rect 269488 57978 269808 58046
rect 269488 57922 269558 57978
rect 269614 57922 269682 57978
rect 269738 57922 269808 57978
rect 269488 57888 269808 57922
rect 300208 58350 300528 58384
rect 300208 58294 300278 58350
rect 300334 58294 300402 58350
rect 300458 58294 300528 58350
rect 300208 58226 300528 58294
rect 300208 58170 300278 58226
rect 300334 58170 300402 58226
rect 300458 58170 300528 58226
rect 300208 58102 300528 58170
rect 300208 58046 300278 58102
rect 300334 58046 300402 58102
rect 300458 58046 300528 58102
rect 300208 57978 300528 58046
rect 300208 57922 300278 57978
rect 300334 57922 300402 57978
rect 300458 57922 300528 57978
rect 300208 57888 300528 57922
rect 330928 58350 331248 58384
rect 330928 58294 330998 58350
rect 331054 58294 331122 58350
rect 331178 58294 331248 58350
rect 330928 58226 331248 58294
rect 330928 58170 330998 58226
rect 331054 58170 331122 58226
rect 331178 58170 331248 58226
rect 330928 58102 331248 58170
rect 330928 58046 330998 58102
rect 331054 58046 331122 58102
rect 331178 58046 331248 58102
rect 330928 57978 331248 58046
rect 330928 57922 330998 57978
rect 331054 57922 331122 57978
rect 331178 57922 331248 57978
rect 330928 57888 331248 57922
rect 361648 58350 361968 58384
rect 361648 58294 361718 58350
rect 361774 58294 361842 58350
rect 361898 58294 361968 58350
rect 361648 58226 361968 58294
rect 361648 58170 361718 58226
rect 361774 58170 361842 58226
rect 361898 58170 361968 58226
rect 361648 58102 361968 58170
rect 361648 58046 361718 58102
rect 361774 58046 361842 58102
rect 361898 58046 361968 58102
rect 361648 57978 361968 58046
rect 361648 57922 361718 57978
rect 361774 57922 361842 57978
rect 361898 57922 361968 57978
rect 361648 57888 361968 57922
rect 392368 58350 392688 58384
rect 392368 58294 392438 58350
rect 392494 58294 392562 58350
rect 392618 58294 392688 58350
rect 392368 58226 392688 58294
rect 392368 58170 392438 58226
rect 392494 58170 392562 58226
rect 392618 58170 392688 58226
rect 392368 58102 392688 58170
rect 392368 58046 392438 58102
rect 392494 58046 392562 58102
rect 392618 58046 392688 58102
rect 392368 57978 392688 58046
rect 392368 57922 392438 57978
rect 392494 57922 392562 57978
rect 392618 57922 392688 57978
rect 392368 57888 392688 57922
rect 423088 58350 423408 58384
rect 423088 58294 423158 58350
rect 423214 58294 423282 58350
rect 423338 58294 423408 58350
rect 423088 58226 423408 58294
rect 423088 58170 423158 58226
rect 423214 58170 423282 58226
rect 423338 58170 423408 58226
rect 423088 58102 423408 58170
rect 423088 58046 423158 58102
rect 423214 58046 423282 58102
rect 423338 58046 423408 58102
rect 423088 57978 423408 58046
rect 423088 57922 423158 57978
rect 423214 57922 423282 57978
rect 423338 57922 423408 57978
rect 423088 57888 423408 57922
rect 453808 58350 454128 58384
rect 453808 58294 453878 58350
rect 453934 58294 454002 58350
rect 454058 58294 454128 58350
rect 453808 58226 454128 58294
rect 453808 58170 453878 58226
rect 453934 58170 454002 58226
rect 454058 58170 454128 58226
rect 453808 58102 454128 58170
rect 453808 58046 453878 58102
rect 453934 58046 454002 58102
rect 454058 58046 454128 58102
rect 453808 57978 454128 58046
rect 453808 57922 453878 57978
rect 453934 57922 454002 57978
rect 454058 57922 454128 57978
rect 453808 57888 454128 57922
rect 484528 58350 484848 58384
rect 484528 58294 484598 58350
rect 484654 58294 484722 58350
rect 484778 58294 484848 58350
rect 484528 58226 484848 58294
rect 484528 58170 484598 58226
rect 484654 58170 484722 58226
rect 484778 58170 484848 58226
rect 484528 58102 484848 58170
rect 484528 58046 484598 58102
rect 484654 58046 484722 58102
rect 484778 58046 484848 58102
rect 484528 57978 484848 58046
rect 484528 57922 484598 57978
rect 484654 57922 484722 57978
rect 484778 57922 484848 57978
rect 484528 57888 484848 57922
rect 515248 58350 515568 58384
rect 515248 58294 515318 58350
rect 515374 58294 515442 58350
rect 515498 58294 515568 58350
rect 515248 58226 515568 58294
rect 515248 58170 515318 58226
rect 515374 58170 515442 58226
rect 515498 58170 515568 58226
rect 515248 58102 515568 58170
rect 515248 58046 515318 58102
rect 515374 58046 515442 58102
rect 515498 58046 515568 58102
rect 515248 57978 515568 58046
rect 515248 57922 515318 57978
rect 515374 57922 515442 57978
rect 515498 57922 515568 57978
rect 515248 57888 515568 57922
rect 545968 58350 546288 58384
rect 545968 58294 546038 58350
rect 546094 58294 546162 58350
rect 546218 58294 546288 58350
rect 545968 58226 546288 58294
rect 545968 58170 546038 58226
rect 546094 58170 546162 58226
rect 546218 58170 546288 58226
rect 545968 58102 546288 58170
rect 545968 58046 546038 58102
rect 546094 58046 546162 58102
rect 546218 58046 546288 58102
rect 545968 57978 546288 58046
rect 545968 57922 546038 57978
rect 546094 57922 546162 57978
rect 546218 57922 546288 57978
rect 545968 57888 546288 57922
rect 561154 58350 561774 75922
rect 561154 58294 561250 58350
rect 561306 58294 561374 58350
rect 561430 58294 561498 58350
rect 561554 58294 561622 58350
rect 561678 58294 561774 58350
rect 561154 58226 561774 58294
rect 561154 58170 561250 58226
rect 561306 58170 561374 58226
rect 561430 58170 561498 58226
rect 561554 58170 561622 58226
rect 561678 58170 561774 58226
rect 561154 58102 561774 58170
rect 561154 58046 561250 58102
rect 561306 58046 561374 58102
rect 561430 58046 561498 58102
rect 561554 58046 561622 58102
rect 561678 58046 561774 58102
rect 561154 57978 561774 58046
rect 561154 57922 561250 57978
rect 561306 57922 561374 57978
rect 561430 57922 561498 57978
rect 561554 57922 561622 57978
rect 561678 57922 561774 57978
rect 131248 46350 131568 46384
rect 131248 46294 131318 46350
rect 131374 46294 131442 46350
rect 131498 46294 131568 46350
rect 131248 46226 131568 46294
rect 131248 46170 131318 46226
rect 131374 46170 131442 46226
rect 131498 46170 131568 46226
rect 131248 46102 131568 46170
rect 131248 46046 131318 46102
rect 131374 46046 131442 46102
rect 131498 46046 131568 46102
rect 131248 45978 131568 46046
rect 131248 45922 131318 45978
rect 131374 45922 131442 45978
rect 131498 45922 131568 45978
rect 131248 45888 131568 45922
rect 161968 46350 162288 46384
rect 161968 46294 162038 46350
rect 162094 46294 162162 46350
rect 162218 46294 162288 46350
rect 161968 46226 162288 46294
rect 161968 46170 162038 46226
rect 162094 46170 162162 46226
rect 162218 46170 162288 46226
rect 161968 46102 162288 46170
rect 161968 46046 162038 46102
rect 162094 46046 162162 46102
rect 162218 46046 162288 46102
rect 161968 45978 162288 46046
rect 161968 45922 162038 45978
rect 162094 45922 162162 45978
rect 162218 45922 162288 45978
rect 161968 45888 162288 45922
rect 192688 46350 193008 46384
rect 192688 46294 192758 46350
rect 192814 46294 192882 46350
rect 192938 46294 193008 46350
rect 192688 46226 193008 46294
rect 192688 46170 192758 46226
rect 192814 46170 192882 46226
rect 192938 46170 193008 46226
rect 192688 46102 193008 46170
rect 192688 46046 192758 46102
rect 192814 46046 192882 46102
rect 192938 46046 193008 46102
rect 192688 45978 193008 46046
rect 192688 45922 192758 45978
rect 192814 45922 192882 45978
rect 192938 45922 193008 45978
rect 192688 45888 193008 45922
rect 223408 46350 223728 46384
rect 223408 46294 223478 46350
rect 223534 46294 223602 46350
rect 223658 46294 223728 46350
rect 223408 46226 223728 46294
rect 223408 46170 223478 46226
rect 223534 46170 223602 46226
rect 223658 46170 223728 46226
rect 223408 46102 223728 46170
rect 223408 46046 223478 46102
rect 223534 46046 223602 46102
rect 223658 46046 223728 46102
rect 223408 45978 223728 46046
rect 223408 45922 223478 45978
rect 223534 45922 223602 45978
rect 223658 45922 223728 45978
rect 223408 45888 223728 45922
rect 254128 46350 254448 46384
rect 254128 46294 254198 46350
rect 254254 46294 254322 46350
rect 254378 46294 254448 46350
rect 254128 46226 254448 46294
rect 254128 46170 254198 46226
rect 254254 46170 254322 46226
rect 254378 46170 254448 46226
rect 254128 46102 254448 46170
rect 254128 46046 254198 46102
rect 254254 46046 254322 46102
rect 254378 46046 254448 46102
rect 254128 45978 254448 46046
rect 254128 45922 254198 45978
rect 254254 45922 254322 45978
rect 254378 45922 254448 45978
rect 254128 45888 254448 45922
rect 284848 46350 285168 46384
rect 284848 46294 284918 46350
rect 284974 46294 285042 46350
rect 285098 46294 285168 46350
rect 284848 46226 285168 46294
rect 284848 46170 284918 46226
rect 284974 46170 285042 46226
rect 285098 46170 285168 46226
rect 284848 46102 285168 46170
rect 284848 46046 284918 46102
rect 284974 46046 285042 46102
rect 285098 46046 285168 46102
rect 284848 45978 285168 46046
rect 284848 45922 284918 45978
rect 284974 45922 285042 45978
rect 285098 45922 285168 45978
rect 284848 45888 285168 45922
rect 315568 46350 315888 46384
rect 315568 46294 315638 46350
rect 315694 46294 315762 46350
rect 315818 46294 315888 46350
rect 315568 46226 315888 46294
rect 315568 46170 315638 46226
rect 315694 46170 315762 46226
rect 315818 46170 315888 46226
rect 315568 46102 315888 46170
rect 315568 46046 315638 46102
rect 315694 46046 315762 46102
rect 315818 46046 315888 46102
rect 315568 45978 315888 46046
rect 315568 45922 315638 45978
rect 315694 45922 315762 45978
rect 315818 45922 315888 45978
rect 315568 45888 315888 45922
rect 346288 46350 346608 46384
rect 346288 46294 346358 46350
rect 346414 46294 346482 46350
rect 346538 46294 346608 46350
rect 346288 46226 346608 46294
rect 346288 46170 346358 46226
rect 346414 46170 346482 46226
rect 346538 46170 346608 46226
rect 346288 46102 346608 46170
rect 346288 46046 346358 46102
rect 346414 46046 346482 46102
rect 346538 46046 346608 46102
rect 346288 45978 346608 46046
rect 346288 45922 346358 45978
rect 346414 45922 346482 45978
rect 346538 45922 346608 45978
rect 346288 45888 346608 45922
rect 377008 46350 377328 46384
rect 377008 46294 377078 46350
rect 377134 46294 377202 46350
rect 377258 46294 377328 46350
rect 377008 46226 377328 46294
rect 377008 46170 377078 46226
rect 377134 46170 377202 46226
rect 377258 46170 377328 46226
rect 377008 46102 377328 46170
rect 377008 46046 377078 46102
rect 377134 46046 377202 46102
rect 377258 46046 377328 46102
rect 377008 45978 377328 46046
rect 377008 45922 377078 45978
rect 377134 45922 377202 45978
rect 377258 45922 377328 45978
rect 377008 45888 377328 45922
rect 407728 46350 408048 46384
rect 407728 46294 407798 46350
rect 407854 46294 407922 46350
rect 407978 46294 408048 46350
rect 407728 46226 408048 46294
rect 407728 46170 407798 46226
rect 407854 46170 407922 46226
rect 407978 46170 408048 46226
rect 407728 46102 408048 46170
rect 407728 46046 407798 46102
rect 407854 46046 407922 46102
rect 407978 46046 408048 46102
rect 407728 45978 408048 46046
rect 407728 45922 407798 45978
rect 407854 45922 407922 45978
rect 407978 45922 408048 45978
rect 407728 45888 408048 45922
rect 438448 46350 438768 46384
rect 438448 46294 438518 46350
rect 438574 46294 438642 46350
rect 438698 46294 438768 46350
rect 438448 46226 438768 46294
rect 438448 46170 438518 46226
rect 438574 46170 438642 46226
rect 438698 46170 438768 46226
rect 438448 46102 438768 46170
rect 438448 46046 438518 46102
rect 438574 46046 438642 46102
rect 438698 46046 438768 46102
rect 438448 45978 438768 46046
rect 438448 45922 438518 45978
rect 438574 45922 438642 45978
rect 438698 45922 438768 45978
rect 438448 45888 438768 45922
rect 469168 46350 469488 46384
rect 469168 46294 469238 46350
rect 469294 46294 469362 46350
rect 469418 46294 469488 46350
rect 469168 46226 469488 46294
rect 469168 46170 469238 46226
rect 469294 46170 469362 46226
rect 469418 46170 469488 46226
rect 469168 46102 469488 46170
rect 469168 46046 469238 46102
rect 469294 46046 469362 46102
rect 469418 46046 469488 46102
rect 469168 45978 469488 46046
rect 469168 45922 469238 45978
rect 469294 45922 469362 45978
rect 469418 45922 469488 45978
rect 469168 45888 469488 45922
rect 499888 46350 500208 46384
rect 499888 46294 499958 46350
rect 500014 46294 500082 46350
rect 500138 46294 500208 46350
rect 499888 46226 500208 46294
rect 499888 46170 499958 46226
rect 500014 46170 500082 46226
rect 500138 46170 500208 46226
rect 499888 46102 500208 46170
rect 499888 46046 499958 46102
rect 500014 46046 500082 46102
rect 500138 46046 500208 46102
rect 499888 45978 500208 46046
rect 499888 45922 499958 45978
rect 500014 45922 500082 45978
rect 500138 45922 500208 45978
rect 499888 45888 500208 45922
rect 530608 46350 530928 46384
rect 530608 46294 530678 46350
rect 530734 46294 530802 46350
rect 530858 46294 530928 46350
rect 530608 46226 530928 46294
rect 530608 46170 530678 46226
rect 530734 46170 530802 46226
rect 530858 46170 530928 46226
rect 530608 46102 530928 46170
rect 530608 46046 530678 46102
rect 530734 46046 530802 46102
rect 530858 46046 530928 46102
rect 530608 45978 530928 46046
rect 530608 45922 530678 45978
rect 530734 45922 530802 45978
rect 530858 45922 530928 45978
rect 530608 45888 530928 45922
rect 111154 40294 111250 40350
rect 111306 40294 111374 40350
rect 111430 40294 111498 40350
rect 111554 40294 111622 40350
rect 111678 40294 111774 40350
rect 111154 40226 111774 40294
rect 111154 40170 111250 40226
rect 111306 40170 111374 40226
rect 111430 40170 111498 40226
rect 111554 40170 111622 40226
rect 111678 40170 111774 40226
rect 111154 40102 111774 40170
rect 111154 40046 111250 40102
rect 111306 40046 111374 40102
rect 111430 40046 111498 40102
rect 111554 40046 111622 40102
rect 111678 40046 111774 40102
rect 111154 39978 111774 40046
rect 111154 39922 111250 39978
rect 111306 39922 111374 39978
rect 111430 39922 111498 39978
rect 111554 39922 111622 39978
rect 111678 39922 111774 39978
rect 111154 22350 111774 39922
rect 115888 40350 116208 40384
rect 115888 40294 115958 40350
rect 116014 40294 116082 40350
rect 116138 40294 116208 40350
rect 115888 40226 116208 40294
rect 115888 40170 115958 40226
rect 116014 40170 116082 40226
rect 116138 40170 116208 40226
rect 115888 40102 116208 40170
rect 115888 40046 115958 40102
rect 116014 40046 116082 40102
rect 116138 40046 116208 40102
rect 115888 39978 116208 40046
rect 115888 39922 115958 39978
rect 116014 39922 116082 39978
rect 116138 39922 116208 39978
rect 115888 39888 116208 39922
rect 146608 40350 146928 40384
rect 146608 40294 146678 40350
rect 146734 40294 146802 40350
rect 146858 40294 146928 40350
rect 146608 40226 146928 40294
rect 146608 40170 146678 40226
rect 146734 40170 146802 40226
rect 146858 40170 146928 40226
rect 146608 40102 146928 40170
rect 146608 40046 146678 40102
rect 146734 40046 146802 40102
rect 146858 40046 146928 40102
rect 146608 39978 146928 40046
rect 146608 39922 146678 39978
rect 146734 39922 146802 39978
rect 146858 39922 146928 39978
rect 146608 39888 146928 39922
rect 177328 40350 177648 40384
rect 177328 40294 177398 40350
rect 177454 40294 177522 40350
rect 177578 40294 177648 40350
rect 177328 40226 177648 40294
rect 177328 40170 177398 40226
rect 177454 40170 177522 40226
rect 177578 40170 177648 40226
rect 177328 40102 177648 40170
rect 177328 40046 177398 40102
rect 177454 40046 177522 40102
rect 177578 40046 177648 40102
rect 177328 39978 177648 40046
rect 177328 39922 177398 39978
rect 177454 39922 177522 39978
rect 177578 39922 177648 39978
rect 177328 39888 177648 39922
rect 208048 40350 208368 40384
rect 208048 40294 208118 40350
rect 208174 40294 208242 40350
rect 208298 40294 208368 40350
rect 208048 40226 208368 40294
rect 208048 40170 208118 40226
rect 208174 40170 208242 40226
rect 208298 40170 208368 40226
rect 208048 40102 208368 40170
rect 208048 40046 208118 40102
rect 208174 40046 208242 40102
rect 208298 40046 208368 40102
rect 208048 39978 208368 40046
rect 208048 39922 208118 39978
rect 208174 39922 208242 39978
rect 208298 39922 208368 39978
rect 208048 39888 208368 39922
rect 238768 40350 239088 40384
rect 238768 40294 238838 40350
rect 238894 40294 238962 40350
rect 239018 40294 239088 40350
rect 238768 40226 239088 40294
rect 238768 40170 238838 40226
rect 238894 40170 238962 40226
rect 239018 40170 239088 40226
rect 238768 40102 239088 40170
rect 238768 40046 238838 40102
rect 238894 40046 238962 40102
rect 239018 40046 239088 40102
rect 238768 39978 239088 40046
rect 238768 39922 238838 39978
rect 238894 39922 238962 39978
rect 239018 39922 239088 39978
rect 238768 39888 239088 39922
rect 269488 40350 269808 40384
rect 269488 40294 269558 40350
rect 269614 40294 269682 40350
rect 269738 40294 269808 40350
rect 269488 40226 269808 40294
rect 269488 40170 269558 40226
rect 269614 40170 269682 40226
rect 269738 40170 269808 40226
rect 269488 40102 269808 40170
rect 269488 40046 269558 40102
rect 269614 40046 269682 40102
rect 269738 40046 269808 40102
rect 269488 39978 269808 40046
rect 269488 39922 269558 39978
rect 269614 39922 269682 39978
rect 269738 39922 269808 39978
rect 269488 39888 269808 39922
rect 300208 40350 300528 40384
rect 300208 40294 300278 40350
rect 300334 40294 300402 40350
rect 300458 40294 300528 40350
rect 300208 40226 300528 40294
rect 300208 40170 300278 40226
rect 300334 40170 300402 40226
rect 300458 40170 300528 40226
rect 300208 40102 300528 40170
rect 300208 40046 300278 40102
rect 300334 40046 300402 40102
rect 300458 40046 300528 40102
rect 300208 39978 300528 40046
rect 300208 39922 300278 39978
rect 300334 39922 300402 39978
rect 300458 39922 300528 39978
rect 300208 39888 300528 39922
rect 330928 40350 331248 40384
rect 330928 40294 330998 40350
rect 331054 40294 331122 40350
rect 331178 40294 331248 40350
rect 330928 40226 331248 40294
rect 330928 40170 330998 40226
rect 331054 40170 331122 40226
rect 331178 40170 331248 40226
rect 330928 40102 331248 40170
rect 330928 40046 330998 40102
rect 331054 40046 331122 40102
rect 331178 40046 331248 40102
rect 330928 39978 331248 40046
rect 330928 39922 330998 39978
rect 331054 39922 331122 39978
rect 331178 39922 331248 39978
rect 330928 39888 331248 39922
rect 361648 40350 361968 40384
rect 361648 40294 361718 40350
rect 361774 40294 361842 40350
rect 361898 40294 361968 40350
rect 361648 40226 361968 40294
rect 361648 40170 361718 40226
rect 361774 40170 361842 40226
rect 361898 40170 361968 40226
rect 361648 40102 361968 40170
rect 361648 40046 361718 40102
rect 361774 40046 361842 40102
rect 361898 40046 361968 40102
rect 361648 39978 361968 40046
rect 361648 39922 361718 39978
rect 361774 39922 361842 39978
rect 361898 39922 361968 39978
rect 361648 39888 361968 39922
rect 392368 40350 392688 40384
rect 392368 40294 392438 40350
rect 392494 40294 392562 40350
rect 392618 40294 392688 40350
rect 392368 40226 392688 40294
rect 392368 40170 392438 40226
rect 392494 40170 392562 40226
rect 392618 40170 392688 40226
rect 392368 40102 392688 40170
rect 392368 40046 392438 40102
rect 392494 40046 392562 40102
rect 392618 40046 392688 40102
rect 392368 39978 392688 40046
rect 392368 39922 392438 39978
rect 392494 39922 392562 39978
rect 392618 39922 392688 39978
rect 392368 39888 392688 39922
rect 423088 40350 423408 40384
rect 423088 40294 423158 40350
rect 423214 40294 423282 40350
rect 423338 40294 423408 40350
rect 423088 40226 423408 40294
rect 423088 40170 423158 40226
rect 423214 40170 423282 40226
rect 423338 40170 423408 40226
rect 423088 40102 423408 40170
rect 423088 40046 423158 40102
rect 423214 40046 423282 40102
rect 423338 40046 423408 40102
rect 423088 39978 423408 40046
rect 423088 39922 423158 39978
rect 423214 39922 423282 39978
rect 423338 39922 423408 39978
rect 423088 39888 423408 39922
rect 453808 40350 454128 40384
rect 453808 40294 453878 40350
rect 453934 40294 454002 40350
rect 454058 40294 454128 40350
rect 453808 40226 454128 40294
rect 453808 40170 453878 40226
rect 453934 40170 454002 40226
rect 454058 40170 454128 40226
rect 453808 40102 454128 40170
rect 453808 40046 453878 40102
rect 453934 40046 454002 40102
rect 454058 40046 454128 40102
rect 453808 39978 454128 40046
rect 453808 39922 453878 39978
rect 453934 39922 454002 39978
rect 454058 39922 454128 39978
rect 453808 39888 454128 39922
rect 484528 40350 484848 40384
rect 484528 40294 484598 40350
rect 484654 40294 484722 40350
rect 484778 40294 484848 40350
rect 484528 40226 484848 40294
rect 484528 40170 484598 40226
rect 484654 40170 484722 40226
rect 484778 40170 484848 40226
rect 484528 40102 484848 40170
rect 484528 40046 484598 40102
rect 484654 40046 484722 40102
rect 484778 40046 484848 40102
rect 484528 39978 484848 40046
rect 484528 39922 484598 39978
rect 484654 39922 484722 39978
rect 484778 39922 484848 39978
rect 484528 39888 484848 39922
rect 515248 40350 515568 40384
rect 515248 40294 515318 40350
rect 515374 40294 515442 40350
rect 515498 40294 515568 40350
rect 515248 40226 515568 40294
rect 515248 40170 515318 40226
rect 515374 40170 515442 40226
rect 515498 40170 515568 40226
rect 515248 40102 515568 40170
rect 515248 40046 515318 40102
rect 515374 40046 515442 40102
rect 515498 40046 515568 40102
rect 515248 39978 515568 40046
rect 515248 39922 515318 39978
rect 515374 39922 515442 39978
rect 515498 39922 515568 39978
rect 515248 39888 515568 39922
rect 545968 40350 546288 40384
rect 545968 40294 546038 40350
rect 546094 40294 546162 40350
rect 546218 40294 546288 40350
rect 545968 40226 546288 40294
rect 545968 40170 546038 40226
rect 546094 40170 546162 40226
rect 546218 40170 546288 40226
rect 545968 40102 546288 40170
rect 545968 40046 546038 40102
rect 546094 40046 546162 40102
rect 546218 40046 546288 40102
rect 545968 39978 546288 40046
rect 545968 39922 546038 39978
rect 546094 39922 546162 39978
rect 546218 39922 546288 39978
rect 545968 39888 546288 39922
rect 561154 40350 561774 57922
rect 561154 40294 561250 40350
rect 561306 40294 561374 40350
rect 561430 40294 561498 40350
rect 561554 40294 561622 40350
rect 561678 40294 561774 40350
rect 561154 40226 561774 40294
rect 561154 40170 561250 40226
rect 561306 40170 561374 40226
rect 561430 40170 561498 40226
rect 561554 40170 561622 40226
rect 561678 40170 561774 40226
rect 561154 40102 561774 40170
rect 561154 40046 561250 40102
rect 561306 40046 561374 40102
rect 561430 40046 561498 40102
rect 561554 40046 561622 40102
rect 561678 40046 561774 40102
rect 561154 39978 561774 40046
rect 561154 39922 561250 39978
rect 561306 39922 561374 39978
rect 561430 39922 561498 39978
rect 561554 39922 561622 39978
rect 561678 39922 561774 39978
rect 111154 22294 111250 22350
rect 111306 22294 111374 22350
rect 111430 22294 111498 22350
rect 111554 22294 111622 22350
rect 111678 22294 111774 22350
rect 111154 22226 111774 22294
rect 111154 22170 111250 22226
rect 111306 22170 111374 22226
rect 111430 22170 111498 22226
rect 111554 22170 111622 22226
rect 111678 22170 111774 22226
rect 111154 22102 111774 22170
rect 111154 22046 111250 22102
rect 111306 22046 111374 22102
rect 111430 22046 111498 22102
rect 111554 22046 111622 22102
rect 111678 22046 111774 22102
rect 111154 21978 111774 22046
rect 111154 21922 111250 21978
rect 111306 21922 111374 21978
rect 111430 21922 111498 21978
rect 111554 21922 111622 21978
rect 111678 21922 111774 21978
rect 111154 4350 111774 21922
rect 111154 4294 111250 4350
rect 111306 4294 111374 4350
rect 111430 4294 111498 4350
rect 111554 4294 111622 4350
rect 111678 4294 111774 4350
rect 111154 4226 111774 4294
rect 111154 4170 111250 4226
rect 111306 4170 111374 4226
rect 111430 4170 111498 4226
rect 111554 4170 111622 4226
rect 111678 4170 111774 4226
rect 111154 4102 111774 4170
rect 111154 4046 111250 4102
rect 111306 4046 111374 4102
rect 111430 4046 111498 4102
rect 111554 4046 111622 4102
rect 111678 4046 111774 4102
rect 111154 3978 111774 4046
rect 111154 3922 111250 3978
rect 111306 3922 111374 3978
rect 111430 3922 111498 3978
rect 111554 3922 111622 3978
rect 111678 3922 111774 3978
rect 111154 -160 111774 3922
rect 111154 -216 111250 -160
rect 111306 -216 111374 -160
rect 111430 -216 111498 -160
rect 111554 -216 111622 -160
rect 111678 -216 111774 -160
rect 111154 -284 111774 -216
rect 111154 -340 111250 -284
rect 111306 -340 111374 -284
rect 111430 -340 111498 -284
rect 111554 -340 111622 -284
rect 111678 -340 111774 -284
rect 111154 -408 111774 -340
rect 111154 -464 111250 -408
rect 111306 -464 111374 -408
rect 111430 -464 111498 -408
rect 111554 -464 111622 -408
rect 111678 -464 111774 -408
rect 111154 -532 111774 -464
rect 111154 -588 111250 -532
rect 111306 -588 111374 -532
rect 111430 -588 111498 -532
rect 111554 -588 111622 -532
rect 111678 -588 111774 -532
rect 111154 -1644 111774 -588
rect 114874 28350 115494 32890
rect 114874 28294 114970 28350
rect 115026 28294 115094 28350
rect 115150 28294 115218 28350
rect 115274 28294 115342 28350
rect 115398 28294 115494 28350
rect 114874 28226 115494 28294
rect 114874 28170 114970 28226
rect 115026 28170 115094 28226
rect 115150 28170 115218 28226
rect 115274 28170 115342 28226
rect 115398 28170 115494 28226
rect 114874 28102 115494 28170
rect 114874 28046 114970 28102
rect 115026 28046 115094 28102
rect 115150 28046 115218 28102
rect 115274 28046 115342 28102
rect 115398 28046 115494 28102
rect 114874 27978 115494 28046
rect 114874 27922 114970 27978
rect 115026 27922 115094 27978
rect 115150 27922 115218 27978
rect 115274 27922 115342 27978
rect 115398 27922 115494 27978
rect 114874 10350 115494 27922
rect 114874 10294 114970 10350
rect 115026 10294 115094 10350
rect 115150 10294 115218 10350
rect 115274 10294 115342 10350
rect 115398 10294 115494 10350
rect 114874 10226 115494 10294
rect 114874 10170 114970 10226
rect 115026 10170 115094 10226
rect 115150 10170 115218 10226
rect 115274 10170 115342 10226
rect 115398 10170 115494 10226
rect 114874 10102 115494 10170
rect 114874 10046 114970 10102
rect 115026 10046 115094 10102
rect 115150 10046 115218 10102
rect 115274 10046 115342 10102
rect 115398 10046 115494 10102
rect 114874 9978 115494 10046
rect 114874 9922 114970 9978
rect 115026 9922 115094 9978
rect 115150 9922 115218 9978
rect 115274 9922 115342 9978
rect 115398 9922 115494 9978
rect 114874 -1120 115494 9922
rect 114874 -1176 114970 -1120
rect 115026 -1176 115094 -1120
rect 115150 -1176 115218 -1120
rect 115274 -1176 115342 -1120
rect 115398 -1176 115494 -1120
rect 114874 -1244 115494 -1176
rect 114874 -1300 114970 -1244
rect 115026 -1300 115094 -1244
rect 115150 -1300 115218 -1244
rect 115274 -1300 115342 -1244
rect 115398 -1300 115494 -1244
rect 114874 -1368 115494 -1300
rect 114874 -1424 114970 -1368
rect 115026 -1424 115094 -1368
rect 115150 -1424 115218 -1368
rect 115274 -1424 115342 -1368
rect 115398 -1424 115494 -1368
rect 114874 -1492 115494 -1424
rect 114874 -1548 114970 -1492
rect 115026 -1548 115094 -1492
rect 115150 -1548 115218 -1492
rect 115274 -1548 115342 -1492
rect 115398 -1548 115494 -1492
rect 114874 -1644 115494 -1548
rect 129154 22350 129774 32890
rect 129154 22294 129250 22350
rect 129306 22294 129374 22350
rect 129430 22294 129498 22350
rect 129554 22294 129622 22350
rect 129678 22294 129774 22350
rect 129154 22226 129774 22294
rect 129154 22170 129250 22226
rect 129306 22170 129374 22226
rect 129430 22170 129498 22226
rect 129554 22170 129622 22226
rect 129678 22170 129774 22226
rect 129154 22102 129774 22170
rect 129154 22046 129250 22102
rect 129306 22046 129374 22102
rect 129430 22046 129498 22102
rect 129554 22046 129622 22102
rect 129678 22046 129774 22102
rect 129154 21978 129774 22046
rect 129154 21922 129250 21978
rect 129306 21922 129374 21978
rect 129430 21922 129498 21978
rect 129554 21922 129622 21978
rect 129678 21922 129774 21978
rect 129154 4350 129774 21922
rect 129154 4294 129250 4350
rect 129306 4294 129374 4350
rect 129430 4294 129498 4350
rect 129554 4294 129622 4350
rect 129678 4294 129774 4350
rect 129154 4226 129774 4294
rect 129154 4170 129250 4226
rect 129306 4170 129374 4226
rect 129430 4170 129498 4226
rect 129554 4170 129622 4226
rect 129678 4170 129774 4226
rect 129154 4102 129774 4170
rect 129154 4046 129250 4102
rect 129306 4046 129374 4102
rect 129430 4046 129498 4102
rect 129554 4046 129622 4102
rect 129678 4046 129774 4102
rect 129154 3978 129774 4046
rect 129154 3922 129250 3978
rect 129306 3922 129374 3978
rect 129430 3922 129498 3978
rect 129554 3922 129622 3978
rect 129678 3922 129774 3978
rect 129154 -160 129774 3922
rect 129154 -216 129250 -160
rect 129306 -216 129374 -160
rect 129430 -216 129498 -160
rect 129554 -216 129622 -160
rect 129678 -216 129774 -160
rect 129154 -284 129774 -216
rect 129154 -340 129250 -284
rect 129306 -340 129374 -284
rect 129430 -340 129498 -284
rect 129554 -340 129622 -284
rect 129678 -340 129774 -284
rect 129154 -408 129774 -340
rect 129154 -464 129250 -408
rect 129306 -464 129374 -408
rect 129430 -464 129498 -408
rect 129554 -464 129622 -408
rect 129678 -464 129774 -408
rect 129154 -532 129774 -464
rect 129154 -588 129250 -532
rect 129306 -588 129374 -532
rect 129430 -588 129498 -532
rect 129554 -588 129622 -532
rect 129678 -588 129774 -532
rect 129154 -1644 129774 -588
rect 132874 28350 133494 32890
rect 132874 28294 132970 28350
rect 133026 28294 133094 28350
rect 133150 28294 133218 28350
rect 133274 28294 133342 28350
rect 133398 28294 133494 28350
rect 132874 28226 133494 28294
rect 132874 28170 132970 28226
rect 133026 28170 133094 28226
rect 133150 28170 133218 28226
rect 133274 28170 133342 28226
rect 133398 28170 133494 28226
rect 132874 28102 133494 28170
rect 132874 28046 132970 28102
rect 133026 28046 133094 28102
rect 133150 28046 133218 28102
rect 133274 28046 133342 28102
rect 133398 28046 133494 28102
rect 132874 27978 133494 28046
rect 132874 27922 132970 27978
rect 133026 27922 133094 27978
rect 133150 27922 133218 27978
rect 133274 27922 133342 27978
rect 133398 27922 133494 27978
rect 132874 10350 133494 27922
rect 132874 10294 132970 10350
rect 133026 10294 133094 10350
rect 133150 10294 133218 10350
rect 133274 10294 133342 10350
rect 133398 10294 133494 10350
rect 132874 10226 133494 10294
rect 132874 10170 132970 10226
rect 133026 10170 133094 10226
rect 133150 10170 133218 10226
rect 133274 10170 133342 10226
rect 133398 10170 133494 10226
rect 132874 10102 133494 10170
rect 132874 10046 132970 10102
rect 133026 10046 133094 10102
rect 133150 10046 133218 10102
rect 133274 10046 133342 10102
rect 133398 10046 133494 10102
rect 132874 9978 133494 10046
rect 132874 9922 132970 9978
rect 133026 9922 133094 9978
rect 133150 9922 133218 9978
rect 133274 9922 133342 9978
rect 133398 9922 133494 9978
rect 132874 -1120 133494 9922
rect 132874 -1176 132970 -1120
rect 133026 -1176 133094 -1120
rect 133150 -1176 133218 -1120
rect 133274 -1176 133342 -1120
rect 133398 -1176 133494 -1120
rect 132874 -1244 133494 -1176
rect 132874 -1300 132970 -1244
rect 133026 -1300 133094 -1244
rect 133150 -1300 133218 -1244
rect 133274 -1300 133342 -1244
rect 133398 -1300 133494 -1244
rect 132874 -1368 133494 -1300
rect 132874 -1424 132970 -1368
rect 133026 -1424 133094 -1368
rect 133150 -1424 133218 -1368
rect 133274 -1424 133342 -1368
rect 133398 -1424 133494 -1368
rect 132874 -1492 133494 -1424
rect 132874 -1548 132970 -1492
rect 133026 -1548 133094 -1492
rect 133150 -1548 133218 -1492
rect 133274 -1548 133342 -1492
rect 133398 -1548 133494 -1492
rect 132874 -1644 133494 -1548
rect 147154 22350 147774 32890
rect 147154 22294 147250 22350
rect 147306 22294 147374 22350
rect 147430 22294 147498 22350
rect 147554 22294 147622 22350
rect 147678 22294 147774 22350
rect 147154 22226 147774 22294
rect 147154 22170 147250 22226
rect 147306 22170 147374 22226
rect 147430 22170 147498 22226
rect 147554 22170 147622 22226
rect 147678 22170 147774 22226
rect 147154 22102 147774 22170
rect 147154 22046 147250 22102
rect 147306 22046 147374 22102
rect 147430 22046 147498 22102
rect 147554 22046 147622 22102
rect 147678 22046 147774 22102
rect 147154 21978 147774 22046
rect 147154 21922 147250 21978
rect 147306 21922 147374 21978
rect 147430 21922 147498 21978
rect 147554 21922 147622 21978
rect 147678 21922 147774 21978
rect 147154 4350 147774 21922
rect 147154 4294 147250 4350
rect 147306 4294 147374 4350
rect 147430 4294 147498 4350
rect 147554 4294 147622 4350
rect 147678 4294 147774 4350
rect 147154 4226 147774 4294
rect 147154 4170 147250 4226
rect 147306 4170 147374 4226
rect 147430 4170 147498 4226
rect 147554 4170 147622 4226
rect 147678 4170 147774 4226
rect 147154 4102 147774 4170
rect 147154 4046 147250 4102
rect 147306 4046 147374 4102
rect 147430 4046 147498 4102
rect 147554 4046 147622 4102
rect 147678 4046 147774 4102
rect 147154 3978 147774 4046
rect 147154 3922 147250 3978
rect 147306 3922 147374 3978
rect 147430 3922 147498 3978
rect 147554 3922 147622 3978
rect 147678 3922 147774 3978
rect 147154 -160 147774 3922
rect 147154 -216 147250 -160
rect 147306 -216 147374 -160
rect 147430 -216 147498 -160
rect 147554 -216 147622 -160
rect 147678 -216 147774 -160
rect 147154 -284 147774 -216
rect 147154 -340 147250 -284
rect 147306 -340 147374 -284
rect 147430 -340 147498 -284
rect 147554 -340 147622 -284
rect 147678 -340 147774 -284
rect 147154 -408 147774 -340
rect 147154 -464 147250 -408
rect 147306 -464 147374 -408
rect 147430 -464 147498 -408
rect 147554 -464 147622 -408
rect 147678 -464 147774 -408
rect 147154 -532 147774 -464
rect 147154 -588 147250 -532
rect 147306 -588 147374 -532
rect 147430 -588 147498 -532
rect 147554 -588 147622 -532
rect 147678 -588 147774 -532
rect 147154 -1644 147774 -588
rect 150874 28350 151494 32890
rect 150874 28294 150970 28350
rect 151026 28294 151094 28350
rect 151150 28294 151218 28350
rect 151274 28294 151342 28350
rect 151398 28294 151494 28350
rect 150874 28226 151494 28294
rect 150874 28170 150970 28226
rect 151026 28170 151094 28226
rect 151150 28170 151218 28226
rect 151274 28170 151342 28226
rect 151398 28170 151494 28226
rect 150874 28102 151494 28170
rect 150874 28046 150970 28102
rect 151026 28046 151094 28102
rect 151150 28046 151218 28102
rect 151274 28046 151342 28102
rect 151398 28046 151494 28102
rect 150874 27978 151494 28046
rect 150874 27922 150970 27978
rect 151026 27922 151094 27978
rect 151150 27922 151218 27978
rect 151274 27922 151342 27978
rect 151398 27922 151494 27978
rect 150874 10350 151494 27922
rect 150874 10294 150970 10350
rect 151026 10294 151094 10350
rect 151150 10294 151218 10350
rect 151274 10294 151342 10350
rect 151398 10294 151494 10350
rect 150874 10226 151494 10294
rect 150874 10170 150970 10226
rect 151026 10170 151094 10226
rect 151150 10170 151218 10226
rect 151274 10170 151342 10226
rect 151398 10170 151494 10226
rect 150874 10102 151494 10170
rect 150874 10046 150970 10102
rect 151026 10046 151094 10102
rect 151150 10046 151218 10102
rect 151274 10046 151342 10102
rect 151398 10046 151494 10102
rect 150874 9978 151494 10046
rect 150874 9922 150970 9978
rect 151026 9922 151094 9978
rect 151150 9922 151218 9978
rect 151274 9922 151342 9978
rect 151398 9922 151494 9978
rect 150874 -1120 151494 9922
rect 150874 -1176 150970 -1120
rect 151026 -1176 151094 -1120
rect 151150 -1176 151218 -1120
rect 151274 -1176 151342 -1120
rect 151398 -1176 151494 -1120
rect 150874 -1244 151494 -1176
rect 150874 -1300 150970 -1244
rect 151026 -1300 151094 -1244
rect 151150 -1300 151218 -1244
rect 151274 -1300 151342 -1244
rect 151398 -1300 151494 -1244
rect 150874 -1368 151494 -1300
rect 150874 -1424 150970 -1368
rect 151026 -1424 151094 -1368
rect 151150 -1424 151218 -1368
rect 151274 -1424 151342 -1368
rect 151398 -1424 151494 -1368
rect 150874 -1492 151494 -1424
rect 150874 -1548 150970 -1492
rect 151026 -1548 151094 -1492
rect 151150 -1548 151218 -1492
rect 151274 -1548 151342 -1492
rect 151398 -1548 151494 -1492
rect 150874 -1644 151494 -1548
rect 165154 22350 165774 32890
rect 165154 22294 165250 22350
rect 165306 22294 165374 22350
rect 165430 22294 165498 22350
rect 165554 22294 165622 22350
rect 165678 22294 165774 22350
rect 165154 22226 165774 22294
rect 165154 22170 165250 22226
rect 165306 22170 165374 22226
rect 165430 22170 165498 22226
rect 165554 22170 165622 22226
rect 165678 22170 165774 22226
rect 165154 22102 165774 22170
rect 165154 22046 165250 22102
rect 165306 22046 165374 22102
rect 165430 22046 165498 22102
rect 165554 22046 165622 22102
rect 165678 22046 165774 22102
rect 165154 21978 165774 22046
rect 165154 21922 165250 21978
rect 165306 21922 165374 21978
rect 165430 21922 165498 21978
rect 165554 21922 165622 21978
rect 165678 21922 165774 21978
rect 165154 4350 165774 21922
rect 165154 4294 165250 4350
rect 165306 4294 165374 4350
rect 165430 4294 165498 4350
rect 165554 4294 165622 4350
rect 165678 4294 165774 4350
rect 165154 4226 165774 4294
rect 165154 4170 165250 4226
rect 165306 4170 165374 4226
rect 165430 4170 165498 4226
rect 165554 4170 165622 4226
rect 165678 4170 165774 4226
rect 165154 4102 165774 4170
rect 165154 4046 165250 4102
rect 165306 4046 165374 4102
rect 165430 4046 165498 4102
rect 165554 4046 165622 4102
rect 165678 4046 165774 4102
rect 165154 3978 165774 4046
rect 165154 3922 165250 3978
rect 165306 3922 165374 3978
rect 165430 3922 165498 3978
rect 165554 3922 165622 3978
rect 165678 3922 165774 3978
rect 165154 -160 165774 3922
rect 165154 -216 165250 -160
rect 165306 -216 165374 -160
rect 165430 -216 165498 -160
rect 165554 -216 165622 -160
rect 165678 -216 165774 -160
rect 165154 -284 165774 -216
rect 165154 -340 165250 -284
rect 165306 -340 165374 -284
rect 165430 -340 165498 -284
rect 165554 -340 165622 -284
rect 165678 -340 165774 -284
rect 165154 -408 165774 -340
rect 165154 -464 165250 -408
rect 165306 -464 165374 -408
rect 165430 -464 165498 -408
rect 165554 -464 165622 -408
rect 165678 -464 165774 -408
rect 165154 -532 165774 -464
rect 165154 -588 165250 -532
rect 165306 -588 165374 -532
rect 165430 -588 165498 -532
rect 165554 -588 165622 -532
rect 165678 -588 165774 -532
rect 165154 -1644 165774 -588
rect 168874 28350 169494 32890
rect 168874 28294 168970 28350
rect 169026 28294 169094 28350
rect 169150 28294 169218 28350
rect 169274 28294 169342 28350
rect 169398 28294 169494 28350
rect 168874 28226 169494 28294
rect 168874 28170 168970 28226
rect 169026 28170 169094 28226
rect 169150 28170 169218 28226
rect 169274 28170 169342 28226
rect 169398 28170 169494 28226
rect 168874 28102 169494 28170
rect 168874 28046 168970 28102
rect 169026 28046 169094 28102
rect 169150 28046 169218 28102
rect 169274 28046 169342 28102
rect 169398 28046 169494 28102
rect 168874 27978 169494 28046
rect 168874 27922 168970 27978
rect 169026 27922 169094 27978
rect 169150 27922 169218 27978
rect 169274 27922 169342 27978
rect 169398 27922 169494 27978
rect 168874 10350 169494 27922
rect 168874 10294 168970 10350
rect 169026 10294 169094 10350
rect 169150 10294 169218 10350
rect 169274 10294 169342 10350
rect 169398 10294 169494 10350
rect 168874 10226 169494 10294
rect 168874 10170 168970 10226
rect 169026 10170 169094 10226
rect 169150 10170 169218 10226
rect 169274 10170 169342 10226
rect 169398 10170 169494 10226
rect 168874 10102 169494 10170
rect 168874 10046 168970 10102
rect 169026 10046 169094 10102
rect 169150 10046 169218 10102
rect 169274 10046 169342 10102
rect 169398 10046 169494 10102
rect 168874 9978 169494 10046
rect 168874 9922 168970 9978
rect 169026 9922 169094 9978
rect 169150 9922 169218 9978
rect 169274 9922 169342 9978
rect 169398 9922 169494 9978
rect 168874 -1120 169494 9922
rect 168874 -1176 168970 -1120
rect 169026 -1176 169094 -1120
rect 169150 -1176 169218 -1120
rect 169274 -1176 169342 -1120
rect 169398 -1176 169494 -1120
rect 168874 -1244 169494 -1176
rect 168874 -1300 168970 -1244
rect 169026 -1300 169094 -1244
rect 169150 -1300 169218 -1244
rect 169274 -1300 169342 -1244
rect 169398 -1300 169494 -1244
rect 168874 -1368 169494 -1300
rect 168874 -1424 168970 -1368
rect 169026 -1424 169094 -1368
rect 169150 -1424 169218 -1368
rect 169274 -1424 169342 -1368
rect 169398 -1424 169494 -1368
rect 168874 -1492 169494 -1424
rect 168874 -1548 168970 -1492
rect 169026 -1548 169094 -1492
rect 169150 -1548 169218 -1492
rect 169274 -1548 169342 -1492
rect 169398 -1548 169494 -1492
rect 168874 -1644 169494 -1548
rect 183154 22350 183774 32890
rect 183154 22294 183250 22350
rect 183306 22294 183374 22350
rect 183430 22294 183498 22350
rect 183554 22294 183622 22350
rect 183678 22294 183774 22350
rect 183154 22226 183774 22294
rect 183154 22170 183250 22226
rect 183306 22170 183374 22226
rect 183430 22170 183498 22226
rect 183554 22170 183622 22226
rect 183678 22170 183774 22226
rect 183154 22102 183774 22170
rect 183154 22046 183250 22102
rect 183306 22046 183374 22102
rect 183430 22046 183498 22102
rect 183554 22046 183622 22102
rect 183678 22046 183774 22102
rect 183154 21978 183774 22046
rect 183154 21922 183250 21978
rect 183306 21922 183374 21978
rect 183430 21922 183498 21978
rect 183554 21922 183622 21978
rect 183678 21922 183774 21978
rect 183154 4350 183774 21922
rect 183154 4294 183250 4350
rect 183306 4294 183374 4350
rect 183430 4294 183498 4350
rect 183554 4294 183622 4350
rect 183678 4294 183774 4350
rect 183154 4226 183774 4294
rect 183154 4170 183250 4226
rect 183306 4170 183374 4226
rect 183430 4170 183498 4226
rect 183554 4170 183622 4226
rect 183678 4170 183774 4226
rect 183154 4102 183774 4170
rect 183154 4046 183250 4102
rect 183306 4046 183374 4102
rect 183430 4046 183498 4102
rect 183554 4046 183622 4102
rect 183678 4046 183774 4102
rect 183154 3978 183774 4046
rect 183154 3922 183250 3978
rect 183306 3922 183374 3978
rect 183430 3922 183498 3978
rect 183554 3922 183622 3978
rect 183678 3922 183774 3978
rect 183154 -160 183774 3922
rect 183154 -216 183250 -160
rect 183306 -216 183374 -160
rect 183430 -216 183498 -160
rect 183554 -216 183622 -160
rect 183678 -216 183774 -160
rect 183154 -284 183774 -216
rect 183154 -340 183250 -284
rect 183306 -340 183374 -284
rect 183430 -340 183498 -284
rect 183554 -340 183622 -284
rect 183678 -340 183774 -284
rect 183154 -408 183774 -340
rect 183154 -464 183250 -408
rect 183306 -464 183374 -408
rect 183430 -464 183498 -408
rect 183554 -464 183622 -408
rect 183678 -464 183774 -408
rect 183154 -532 183774 -464
rect 183154 -588 183250 -532
rect 183306 -588 183374 -532
rect 183430 -588 183498 -532
rect 183554 -588 183622 -532
rect 183678 -588 183774 -532
rect 183154 -1644 183774 -588
rect 186874 28350 187494 32890
rect 186874 28294 186970 28350
rect 187026 28294 187094 28350
rect 187150 28294 187218 28350
rect 187274 28294 187342 28350
rect 187398 28294 187494 28350
rect 186874 28226 187494 28294
rect 186874 28170 186970 28226
rect 187026 28170 187094 28226
rect 187150 28170 187218 28226
rect 187274 28170 187342 28226
rect 187398 28170 187494 28226
rect 186874 28102 187494 28170
rect 186874 28046 186970 28102
rect 187026 28046 187094 28102
rect 187150 28046 187218 28102
rect 187274 28046 187342 28102
rect 187398 28046 187494 28102
rect 186874 27978 187494 28046
rect 186874 27922 186970 27978
rect 187026 27922 187094 27978
rect 187150 27922 187218 27978
rect 187274 27922 187342 27978
rect 187398 27922 187494 27978
rect 186874 10350 187494 27922
rect 186874 10294 186970 10350
rect 187026 10294 187094 10350
rect 187150 10294 187218 10350
rect 187274 10294 187342 10350
rect 187398 10294 187494 10350
rect 186874 10226 187494 10294
rect 186874 10170 186970 10226
rect 187026 10170 187094 10226
rect 187150 10170 187218 10226
rect 187274 10170 187342 10226
rect 187398 10170 187494 10226
rect 186874 10102 187494 10170
rect 186874 10046 186970 10102
rect 187026 10046 187094 10102
rect 187150 10046 187218 10102
rect 187274 10046 187342 10102
rect 187398 10046 187494 10102
rect 186874 9978 187494 10046
rect 186874 9922 186970 9978
rect 187026 9922 187094 9978
rect 187150 9922 187218 9978
rect 187274 9922 187342 9978
rect 187398 9922 187494 9978
rect 186874 -1120 187494 9922
rect 186874 -1176 186970 -1120
rect 187026 -1176 187094 -1120
rect 187150 -1176 187218 -1120
rect 187274 -1176 187342 -1120
rect 187398 -1176 187494 -1120
rect 186874 -1244 187494 -1176
rect 186874 -1300 186970 -1244
rect 187026 -1300 187094 -1244
rect 187150 -1300 187218 -1244
rect 187274 -1300 187342 -1244
rect 187398 -1300 187494 -1244
rect 186874 -1368 187494 -1300
rect 186874 -1424 186970 -1368
rect 187026 -1424 187094 -1368
rect 187150 -1424 187218 -1368
rect 187274 -1424 187342 -1368
rect 187398 -1424 187494 -1368
rect 186874 -1492 187494 -1424
rect 186874 -1548 186970 -1492
rect 187026 -1548 187094 -1492
rect 187150 -1548 187218 -1492
rect 187274 -1548 187342 -1492
rect 187398 -1548 187494 -1492
rect 186874 -1644 187494 -1548
rect 201154 22350 201774 32890
rect 201154 22294 201250 22350
rect 201306 22294 201374 22350
rect 201430 22294 201498 22350
rect 201554 22294 201622 22350
rect 201678 22294 201774 22350
rect 201154 22226 201774 22294
rect 201154 22170 201250 22226
rect 201306 22170 201374 22226
rect 201430 22170 201498 22226
rect 201554 22170 201622 22226
rect 201678 22170 201774 22226
rect 201154 22102 201774 22170
rect 201154 22046 201250 22102
rect 201306 22046 201374 22102
rect 201430 22046 201498 22102
rect 201554 22046 201622 22102
rect 201678 22046 201774 22102
rect 201154 21978 201774 22046
rect 201154 21922 201250 21978
rect 201306 21922 201374 21978
rect 201430 21922 201498 21978
rect 201554 21922 201622 21978
rect 201678 21922 201774 21978
rect 201154 4350 201774 21922
rect 201154 4294 201250 4350
rect 201306 4294 201374 4350
rect 201430 4294 201498 4350
rect 201554 4294 201622 4350
rect 201678 4294 201774 4350
rect 201154 4226 201774 4294
rect 201154 4170 201250 4226
rect 201306 4170 201374 4226
rect 201430 4170 201498 4226
rect 201554 4170 201622 4226
rect 201678 4170 201774 4226
rect 201154 4102 201774 4170
rect 201154 4046 201250 4102
rect 201306 4046 201374 4102
rect 201430 4046 201498 4102
rect 201554 4046 201622 4102
rect 201678 4046 201774 4102
rect 201154 3978 201774 4046
rect 201154 3922 201250 3978
rect 201306 3922 201374 3978
rect 201430 3922 201498 3978
rect 201554 3922 201622 3978
rect 201678 3922 201774 3978
rect 201154 -160 201774 3922
rect 201154 -216 201250 -160
rect 201306 -216 201374 -160
rect 201430 -216 201498 -160
rect 201554 -216 201622 -160
rect 201678 -216 201774 -160
rect 201154 -284 201774 -216
rect 201154 -340 201250 -284
rect 201306 -340 201374 -284
rect 201430 -340 201498 -284
rect 201554 -340 201622 -284
rect 201678 -340 201774 -284
rect 201154 -408 201774 -340
rect 201154 -464 201250 -408
rect 201306 -464 201374 -408
rect 201430 -464 201498 -408
rect 201554 -464 201622 -408
rect 201678 -464 201774 -408
rect 201154 -532 201774 -464
rect 201154 -588 201250 -532
rect 201306 -588 201374 -532
rect 201430 -588 201498 -532
rect 201554 -588 201622 -532
rect 201678 -588 201774 -532
rect 201154 -1644 201774 -588
rect 204874 28350 205494 32890
rect 204874 28294 204970 28350
rect 205026 28294 205094 28350
rect 205150 28294 205218 28350
rect 205274 28294 205342 28350
rect 205398 28294 205494 28350
rect 204874 28226 205494 28294
rect 204874 28170 204970 28226
rect 205026 28170 205094 28226
rect 205150 28170 205218 28226
rect 205274 28170 205342 28226
rect 205398 28170 205494 28226
rect 204874 28102 205494 28170
rect 204874 28046 204970 28102
rect 205026 28046 205094 28102
rect 205150 28046 205218 28102
rect 205274 28046 205342 28102
rect 205398 28046 205494 28102
rect 204874 27978 205494 28046
rect 204874 27922 204970 27978
rect 205026 27922 205094 27978
rect 205150 27922 205218 27978
rect 205274 27922 205342 27978
rect 205398 27922 205494 27978
rect 204874 10350 205494 27922
rect 204874 10294 204970 10350
rect 205026 10294 205094 10350
rect 205150 10294 205218 10350
rect 205274 10294 205342 10350
rect 205398 10294 205494 10350
rect 204874 10226 205494 10294
rect 204874 10170 204970 10226
rect 205026 10170 205094 10226
rect 205150 10170 205218 10226
rect 205274 10170 205342 10226
rect 205398 10170 205494 10226
rect 204874 10102 205494 10170
rect 204874 10046 204970 10102
rect 205026 10046 205094 10102
rect 205150 10046 205218 10102
rect 205274 10046 205342 10102
rect 205398 10046 205494 10102
rect 204874 9978 205494 10046
rect 204874 9922 204970 9978
rect 205026 9922 205094 9978
rect 205150 9922 205218 9978
rect 205274 9922 205342 9978
rect 205398 9922 205494 9978
rect 204874 -1120 205494 9922
rect 204874 -1176 204970 -1120
rect 205026 -1176 205094 -1120
rect 205150 -1176 205218 -1120
rect 205274 -1176 205342 -1120
rect 205398 -1176 205494 -1120
rect 204874 -1244 205494 -1176
rect 204874 -1300 204970 -1244
rect 205026 -1300 205094 -1244
rect 205150 -1300 205218 -1244
rect 205274 -1300 205342 -1244
rect 205398 -1300 205494 -1244
rect 204874 -1368 205494 -1300
rect 204874 -1424 204970 -1368
rect 205026 -1424 205094 -1368
rect 205150 -1424 205218 -1368
rect 205274 -1424 205342 -1368
rect 205398 -1424 205494 -1368
rect 204874 -1492 205494 -1424
rect 204874 -1548 204970 -1492
rect 205026 -1548 205094 -1492
rect 205150 -1548 205218 -1492
rect 205274 -1548 205342 -1492
rect 205398 -1548 205494 -1492
rect 204874 -1644 205494 -1548
rect 219154 22350 219774 32890
rect 219154 22294 219250 22350
rect 219306 22294 219374 22350
rect 219430 22294 219498 22350
rect 219554 22294 219622 22350
rect 219678 22294 219774 22350
rect 219154 22226 219774 22294
rect 219154 22170 219250 22226
rect 219306 22170 219374 22226
rect 219430 22170 219498 22226
rect 219554 22170 219622 22226
rect 219678 22170 219774 22226
rect 219154 22102 219774 22170
rect 219154 22046 219250 22102
rect 219306 22046 219374 22102
rect 219430 22046 219498 22102
rect 219554 22046 219622 22102
rect 219678 22046 219774 22102
rect 219154 21978 219774 22046
rect 219154 21922 219250 21978
rect 219306 21922 219374 21978
rect 219430 21922 219498 21978
rect 219554 21922 219622 21978
rect 219678 21922 219774 21978
rect 219154 4350 219774 21922
rect 219154 4294 219250 4350
rect 219306 4294 219374 4350
rect 219430 4294 219498 4350
rect 219554 4294 219622 4350
rect 219678 4294 219774 4350
rect 219154 4226 219774 4294
rect 219154 4170 219250 4226
rect 219306 4170 219374 4226
rect 219430 4170 219498 4226
rect 219554 4170 219622 4226
rect 219678 4170 219774 4226
rect 219154 4102 219774 4170
rect 219154 4046 219250 4102
rect 219306 4046 219374 4102
rect 219430 4046 219498 4102
rect 219554 4046 219622 4102
rect 219678 4046 219774 4102
rect 219154 3978 219774 4046
rect 219154 3922 219250 3978
rect 219306 3922 219374 3978
rect 219430 3922 219498 3978
rect 219554 3922 219622 3978
rect 219678 3922 219774 3978
rect 219154 -160 219774 3922
rect 219154 -216 219250 -160
rect 219306 -216 219374 -160
rect 219430 -216 219498 -160
rect 219554 -216 219622 -160
rect 219678 -216 219774 -160
rect 219154 -284 219774 -216
rect 219154 -340 219250 -284
rect 219306 -340 219374 -284
rect 219430 -340 219498 -284
rect 219554 -340 219622 -284
rect 219678 -340 219774 -284
rect 219154 -408 219774 -340
rect 219154 -464 219250 -408
rect 219306 -464 219374 -408
rect 219430 -464 219498 -408
rect 219554 -464 219622 -408
rect 219678 -464 219774 -408
rect 219154 -532 219774 -464
rect 219154 -588 219250 -532
rect 219306 -588 219374 -532
rect 219430 -588 219498 -532
rect 219554 -588 219622 -532
rect 219678 -588 219774 -532
rect 219154 -1644 219774 -588
rect 222874 28350 223494 31020
rect 222874 28294 222970 28350
rect 223026 28294 223094 28350
rect 223150 28294 223218 28350
rect 223274 28294 223342 28350
rect 223398 28294 223494 28350
rect 222874 28226 223494 28294
rect 222874 28170 222970 28226
rect 223026 28170 223094 28226
rect 223150 28170 223218 28226
rect 223274 28170 223342 28226
rect 223398 28170 223494 28226
rect 222874 28102 223494 28170
rect 222874 28046 222970 28102
rect 223026 28046 223094 28102
rect 223150 28046 223218 28102
rect 223274 28046 223342 28102
rect 223398 28046 223494 28102
rect 222874 27978 223494 28046
rect 222874 27922 222970 27978
rect 223026 27922 223094 27978
rect 223150 27922 223218 27978
rect 223274 27922 223342 27978
rect 223398 27922 223494 27978
rect 222874 10350 223494 27922
rect 222874 10294 222970 10350
rect 223026 10294 223094 10350
rect 223150 10294 223218 10350
rect 223274 10294 223342 10350
rect 223398 10294 223494 10350
rect 222874 10226 223494 10294
rect 222874 10170 222970 10226
rect 223026 10170 223094 10226
rect 223150 10170 223218 10226
rect 223274 10170 223342 10226
rect 223398 10170 223494 10226
rect 222874 10102 223494 10170
rect 222874 10046 222970 10102
rect 223026 10046 223094 10102
rect 223150 10046 223218 10102
rect 223274 10046 223342 10102
rect 223398 10046 223494 10102
rect 222874 9978 223494 10046
rect 222874 9922 222970 9978
rect 223026 9922 223094 9978
rect 223150 9922 223218 9978
rect 223274 9922 223342 9978
rect 223398 9922 223494 9978
rect 222874 -1120 223494 9922
rect 222874 -1176 222970 -1120
rect 223026 -1176 223094 -1120
rect 223150 -1176 223218 -1120
rect 223274 -1176 223342 -1120
rect 223398 -1176 223494 -1120
rect 222874 -1244 223494 -1176
rect 222874 -1300 222970 -1244
rect 223026 -1300 223094 -1244
rect 223150 -1300 223218 -1244
rect 223274 -1300 223342 -1244
rect 223398 -1300 223494 -1244
rect 222874 -1368 223494 -1300
rect 222874 -1424 222970 -1368
rect 223026 -1424 223094 -1368
rect 223150 -1424 223218 -1368
rect 223274 -1424 223342 -1368
rect 223398 -1424 223494 -1368
rect 222874 -1492 223494 -1424
rect 222874 -1548 222970 -1492
rect 223026 -1548 223094 -1492
rect 223150 -1548 223218 -1492
rect 223274 -1548 223342 -1492
rect 223398 -1548 223494 -1492
rect 222874 -1644 223494 -1548
rect 237154 22350 237774 32890
rect 237154 22294 237250 22350
rect 237306 22294 237374 22350
rect 237430 22294 237498 22350
rect 237554 22294 237622 22350
rect 237678 22294 237774 22350
rect 237154 22226 237774 22294
rect 237154 22170 237250 22226
rect 237306 22170 237374 22226
rect 237430 22170 237498 22226
rect 237554 22170 237622 22226
rect 237678 22170 237774 22226
rect 237154 22102 237774 22170
rect 237154 22046 237250 22102
rect 237306 22046 237374 22102
rect 237430 22046 237498 22102
rect 237554 22046 237622 22102
rect 237678 22046 237774 22102
rect 237154 21978 237774 22046
rect 237154 21922 237250 21978
rect 237306 21922 237374 21978
rect 237430 21922 237498 21978
rect 237554 21922 237622 21978
rect 237678 21922 237774 21978
rect 237154 4350 237774 21922
rect 237154 4294 237250 4350
rect 237306 4294 237374 4350
rect 237430 4294 237498 4350
rect 237554 4294 237622 4350
rect 237678 4294 237774 4350
rect 237154 4226 237774 4294
rect 237154 4170 237250 4226
rect 237306 4170 237374 4226
rect 237430 4170 237498 4226
rect 237554 4170 237622 4226
rect 237678 4170 237774 4226
rect 237154 4102 237774 4170
rect 237154 4046 237250 4102
rect 237306 4046 237374 4102
rect 237430 4046 237498 4102
rect 237554 4046 237622 4102
rect 237678 4046 237774 4102
rect 237154 3978 237774 4046
rect 237154 3922 237250 3978
rect 237306 3922 237374 3978
rect 237430 3922 237498 3978
rect 237554 3922 237622 3978
rect 237678 3922 237774 3978
rect 237154 -160 237774 3922
rect 237154 -216 237250 -160
rect 237306 -216 237374 -160
rect 237430 -216 237498 -160
rect 237554 -216 237622 -160
rect 237678 -216 237774 -160
rect 237154 -284 237774 -216
rect 237154 -340 237250 -284
rect 237306 -340 237374 -284
rect 237430 -340 237498 -284
rect 237554 -340 237622 -284
rect 237678 -340 237774 -284
rect 237154 -408 237774 -340
rect 237154 -464 237250 -408
rect 237306 -464 237374 -408
rect 237430 -464 237498 -408
rect 237554 -464 237622 -408
rect 237678 -464 237774 -408
rect 237154 -532 237774 -464
rect 237154 -588 237250 -532
rect 237306 -588 237374 -532
rect 237430 -588 237498 -532
rect 237554 -588 237622 -532
rect 237678 -588 237774 -532
rect 237154 -1644 237774 -588
rect 240874 28350 241494 32890
rect 240874 28294 240970 28350
rect 241026 28294 241094 28350
rect 241150 28294 241218 28350
rect 241274 28294 241342 28350
rect 241398 28294 241494 28350
rect 240874 28226 241494 28294
rect 240874 28170 240970 28226
rect 241026 28170 241094 28226
rect 241150 28170 241218 28226
rect 241274 28170 241342 28226
rect 241398 28170 241494 28226
rect 240874 28102 241494 28170
rect 240874 28046 240970 28102
rect 241026 28046 241094 28102
rect 241150 28046 241218 28102
rect 241274 28046 241342 28102
rect 241398 28046 241494 28102
rect 240874 27978 241494 28046
rect 240874 27922 240970 27978
rect 241026 27922 241094 27978
rect 241150 27922 241218 27978
rect 241274 27922 241342 27978
rect 241398 27922 241494 27978
rect 240874 10350 241494 27922
rect 240874 10294 240970 10350
rect 241026 10294 241094 10350
rect 241150 10294 241218 10350
rect 241274 10294 241342 10350
rect 241398 10294 241494 10350
rect 240874 10226 241494 10294
rect 240874 10170 240970 10226
rect 241026 10170 241094 10226
rect 241150 10170 241218 10226
rect 241274 10170 241342 10226
rect 241398 10170 241494 10226
rect 240874 10102 241494 10170
rect 240874 10046 240970 10102
rect 241026 10046 241094 10102
rect 241150 10046 241218 10102
rect 241274 10046 241342 10102
rect 241398 10046 241494 10102
rect 240874 9978 241494 10046
rect 240874 9922 240970 9978
rect 241026 9922 241094 9978
rect 241150 9922 241218 9978
rect 241274 9922 241342 9978
rect 241398 9922 241494 9978
rect 240874 -1120 241494 9922
rect 240874 -1176 240970 -1120
rect 241026 -1176 241094 -1120
rect 241150 -1176 241218 -1120
rect 241274 -1176 241342 -1120
rect 241398 -1176 241494 -1120
rect 240874 -1244 241494 -1176
rect 240874 -1300 240970 -1244
rect 241026 -1300 241094 -1244
rect 241150 -1300 241218 -1244
rect 241274 -1300 241342 -1244
rect 241398 -1300 241494 -1244
rect 240874 -1368 241494 -1300
rect 240874 -1424 240970 -1368
rect 241026 -1424 241094 -1368
rect 241150 -1424 241218 -1368
rect 241274 -1424 241342 -1368
rect 241398 -1424 241494 -1368
rect 240874 -1492 241494 -1424
rect 240874 -1548 240970 -1492
rect 241026 -1548 241094 -1492
rect 241150 -1548 241218 -1492
rect 241274 -1548 241342 -1492
rect 241398 -1548 241494 -1492
rect 240874 -1644 241494 -1548
rect 255154 22350 255774 32890
rect 255154 22294 255250 22350
rect 255306 22294 255374 22350
rect 255430 22294 255498 22350
rect 255554 22294 255622 22350
rect 255678 22294 255774 22350
rect 255154 22226 255774 22294
rect 255154 22170 255250 22226
rect 255306 22170 255374 22226
rect 255430 22170 255498 22226
rect 255554 22170 255622 22226
rect 255678 22170 255774 22226
rect 255154 22102 255774 22170
rect 255154 22046 255250 22102
rect 255306 22046 255374 22102
rect 255430 22046 255498 22102
rect 255554 22046 255622 22102
rect 255678 22046 255774 22102
rect 255154 21978 255774 22046
rect 255154 21922 255250 21978
rect 255306 21922 255374 21978
rect 255430 21922 255498 21978
rect 255554 21922 255622 21978
rect 255678 21922 255774 21978
rect 255154 4350 255774 21922
rect 255154 4294 255250 4350
rect 255306 4294 255374 4350
rect 255430 4294 255498 4350
rect 255554 4294 255622 4350
rect 255678 4294 255774 4350
rect 255154 4226 255774 4294
rect 255154 4170 255250 4226
rect 255306 4170 255374 4226
rect 255430 4170 255498 4226
rect 255554 4170 255622 4226
rect 255678 4170 255774 4226
rect 255154 4102 255774 4170
rect 255154 4046 255250 4102
rect 255306 4046 255374 4102
rect 255430 4046 255498 4102
rect 255554 4046 255622 4102
rect 255678 4046 255774 4102
rect 255154 3978 255774 4046
rect 255154 3922 255250 3978
rect 255306 3922 255374 3978
rect 255430 3922 255498 3978
rect 255554 3922 255622 3978
rect 255678 3922 255774 3978
rect 255154 -160 255774 3922
rect 255154 -216 255250 -160
rect 255306 -216 255374 -160
rect 255430 -216 255498 -160
rect 255554 -216 255622 -160
rect 255678 -216 255774 -160
rect 255154 -284 255774 -216
rect 255154 -340 255250 -284
rect 255306 -340 255374 -284
rect 255430 -340 255498 -284
rect 255554 -340 255622 -284
rect 255678 -340 255774 -284
rect 255154 -408 255774 -340
rect 255154 -464 255250 -408
rect 255306 -464 255374 -408
rect 255430 -464 255498 -408
rect 255554 -464 255622 -408
rect 255678 -464 255774 -408
rect 255154 -532 255774 -464
rect 255154 -588 255250 -532
rect 255306 -588 255374 -532
rect 255430 -588 255498 -532
rect 255554 -588 255622 -532
rect 255678 -588 255774 -532
rect 255154 -1644 255774 -588
rect 258874 28350 259494 32890
rect 258874 28294 258970 28350
rect 259026 28294 259094 28350
rect 259150 28294 259218 28350
rect 259274 28294 259342 28350
rect 259398 28294 259494 28350
rect 258874 28226 259494 28294
rect 258874 28170 258970 28226
rect 259026 28170 259094 28226
rect 259150 28170 259218 28226
rect 259274 28170 259342 28226
rect 259398 28170 259494 28226
rect 258874 28102 259494 28170
rect 258874 28046 258970 28102
rect 259026 28046 259094 28102
rect 259150 28046 259218 28102
rect 259274 28046 259342 28102
rect 259398 28046 259494 28102
rect 258874 27978 259494 28046
rect 258874 27922 258970 27978
rect 259026 27922 259094 27978
rect 259150 27922 259218 27978
rect 259274 27922 259342 27978
rect 259398 27922 259494 27978
rect 258874 10350 259494 27922
rect 258874 10294 258970 10350
rect 259026 10294 259094 10350
rect 259150 10294 259218 10350
rect 259274 10294 259342 10350
rect 259398 10294 259494 10350
rect 258874 10226 259494 10294
rect 258874 10170 258970 10226
rect 259026 10170 259094 10226
rect 259150 10170 259218 10226
rect 259274 10170 259342 10226
rect 259398 10170 259494 10226
rect 258874 10102 259494 10170
rect 258874 10046 258970 10102
rect 259026 10046 259094 10102
rect 259150 10046 259218 10102
rect 259274 10046 259342 10102
rect 259398 10046 259494 10102
rect 258874 9978 259494 10046
rect 258874 9922 258970 9978
rect 259026 9922 259094 9978
rect 259150 9922 259218 9978
rect 259274 9922 259342 9978
rect 259398 9922 259494 9978
rect 258874 -1120 259494 9922
rect 258874 -1176 258970 -1120
rect 259026 -1176 259094 -1120
rect 259150 -1176 259218 -1120
rect 259274 -1176 259342 -1120
rect 259398 -1176 259494 -1120
rect 258874 -1244 259494 -1176
rect 258874 -1300 258970 -1244
rect 259026 -1300 259094 -1244
rect 259150 -1300 259218 -1244
rect 259274 -1300 259342 -1244
rect 259398 -1300 259494 -1244
rect 258874 -1368 259494 -1300
rect 258874 -1424 258970 -1368
rect 259026 -1424 259094 -1368
rect 259150 -1424 259218 -1368
rect 259274 -1424 259342 -1368
rect 259398 -1424 259494 -1368
rect 258874 -1492 259494 -1424
rect 258874 -1548 258970 -1492
rect 259026 -1548 259094 -1492
rect 259150 -1548 259218 -1492
rect 259274 -1548 259342 -1492
rect 259398 -1548 259494 -1492
rect 258874 -1644 259494 -1548
rect 273154 22350 273774 32890
rect 273154 22294 273250 22350
rect 273306 22294 273374 22350
rect 273430 22294 273498 22350
rect 273554 22294 273622 22350
rect 273678 22294 273774 22350
rect 273154 22226 273774 22294
rect 273154 22170 273250 22226
rect 273306 22170 273374 22226
rect 273430 22170 273498 22226
rect 273554 22170 273622 22226
rect 273678 22170 273774 22226
rect 273154 22102 273774 22170
rect 273154 22046 273250 22102
rect 273306 22046 273374 22102
rect 273430 22046 273498 22102
rect 273554 22046 273622 22102
rect 273678 22046 273774 22102
rect 273154 21978 273774 22046
rect 273154 21922 273250 21978
rect 273306 21922 273374 21978
rect 273430 21922 273498 21978
rect 273554 21922 273622 21978
rect 273678 21922 273774 21978
rect 273154 4350 273774 21922
rect 273154 4294 273250 4350
rect 273306 4294 273374 4350
rect 273430 4294 273498 4350
rect 273554 4294 273622 4350
rect 273678 4294 273774 4350
rect 273154 4226 273774 4294
rect 273154 4170 273250 4226
rect 273306 4170 273374 4226
rect 273430 4170 273498 4226
rect 273554 4170 273622 4226
rect 273678 4170 273774 4226
rect 273154 4102 273774 4170
rect 273154 4046 273250 4102
rect 273306 4046 273374 4102
rect 273430 4046 273498 4102
rect 273554 4046 273622 4102
rect 273678 4046 273774 4102
rect 273154 3978 273774 4046
rect 273154 3922 273250 3978
rect 273306 3922 273374 3978
rect 273430 3922 273498 3978
rect 273554 3922 273622 3978
rect 273678 3922 273774 3978
rect 273154 -160 273774 3922
rect 273154 -216 273250 -160
rect 273306 -216 273374 -160
rect 273430 -216 273498 -160
rect 273554 -216 273622 -160
rect 273678 -216 273774 -160
rect 273154 -284 273774 -216
rect 273154 -340 273250 -284
rect 273306 -340 273374 -284
rect 273430 -340 273498 -284
rect 273554 -340 273622 -284
rect 273678 -340 273774 -284
rect 273154 -408 273774 -340
rect 273154 -464 273250 -408
rect 273306 -464 273374 -408
rect 273430 -464 273498 -408
rect 273554 -464 273622 -408
rect 273678 -464 273774 -408
rect 273154 -532 273774 -464
rect 273154 -588 273250 -532
rect 273306 -588 273374 -532
rect 273430 -588 273498 -532
rect 273554 -588 273622 -532
rect 273678 -588 273774 -532
rect 273154 -1644 273774 -588
rect 276874 28350 277494 32890
rect 276874 28294 276970 28350
rect 277026 28294 277094 28350
rect 277150 28294 277218 28350
rect 277274 28294 277342 28350
rect 277398 28294 277494 28350
rect 276874 28226 277494 28294
rect 276874 28170 276970 28226
rect 277026 28170 277094 28226
rect 277150 28170 277218 28226
rect 277274 28170 277342 28226
rect 277398 28170 277494 28226
rect 276874 28102 277494 28170
rect 276874 28046 276970 28102
rect 277026 28046 277094 28102
rect 277150 28046 277218 28102
rect 277274 28046 277342 28102
rect 277398 28046 277494 28102
rect 276874 27978 277494 28046
rect 276874 27922 276970 27978
rect 277026 27922 277094 27978
rect 277150 27922 277218 27978
rect 277274 27922 277342 27978
rect 277398 27922 277494 27978
rect 276874 10350 277494 27922
rect 276874 10294 276970 10350
rect 277026 10294 277094 10350
rect 277150 10294 277218 10350
rect 277274 10294 277342 10350
rect 277398 10294 277494 10350
rect 276874 10226 277494 10294
rect 276874 10170 276970 10226
rect 277026 10170 277094 10226
rect 277150 10170 277218 10226
rect 277274 10170 277342 10226
rect 277398 10170 277494 10226
rect 276874 10102 277494 10170
rect 276874 10046 276970 10102
rect 277026 10046 277094 10102
rect 277150 10046 277218 10102
rect 277274 10046 277342 10102
rect 277398 10046 277494 10102
rect 276874 9978 277494 10046
rect 276874 9922 276970 9978
rect 277026 9922 277094 9978
rect 277150 9922 277218 9978
rect 277274 9922 277342 9978
rect 277398 9922 277494 9978
rect 276874 -1120 277494 9922
rect 276874 -1176 276970 -1120
rect 277026 -1176 277094 -1120
rect 277150 -1176 277218 -1120
rect 277274 -1176 277342 -1120
rect 277398 -1176 277494 -1120
rect 276874 -1244 277494 -1176
rect 276874 -1300 276970 -1244
rect 277026 -1300 277094 -1244
rect 277150 -1300 277218 -1244
rect 277274 -1300 277342 -1244
rect 277398 -1300 277494 -1244
rect 276874 -1368 277494 -1300
rect 276874 -1424 276970 -1368
rect 277026 -1424 277094 -1368
rect 277150 -1424 277218 -1368
rect 277274 -1424 277342 -1368
rect 277398 -1424 277494 -1368
rect 276874 -1492 277494 -1424
rect 276874 -1548 276970 -1492
rect 277026 -1548 277094 -1492
rect 277150 -1548 277218 -1492
rect 277274 -1548 277342 -1492
rect 277398 -1548 277494 -1492
rect 276874 -1644 277494 -1548
rect 291154 22350 291774 32890
rect 291154 22294 291250 22350
rect 291306 22294 291374 22350
rect 291430 22294 291498 22350
rect 291554 22294 291622 22350
rect 291678 22294 291774 22350
rect 291154 22226 291774 22294
rect 291154 22170 291250 22226
rect 291306 22170 291374 22226
rect 291430 22170 291498 22226
rect 291554 22170 291622 22226
rect 291678 22170 291774 22226
rect 291154 22102 291774 22170
rect 291154 22046 291250 22102
rect 291306 22046 291374 22102
rect 291430 22046 291498 22102
rect 291554 22046 291622 22102
rect 291678 22046 291774 22102
rect 291154 21978 291774 22046
rect 291154 21922 291250 21978
rect 291306 21922 291374 21978
rect 291430 21922 291498 21978
rect 291554 21922 291622 21978
rect 291678 21922 291774 21978
rect 291154 4350 291774 21922
rect 291154 4294 291250 4350
rect 291306 4294 291374 4350
rect 291430 4294 291498 4350
rect 291554 4294 291622 4350
rect 291678 4294 291774 4350
rect 291154 4226 291774 4294
rect 291154 4170 291250 4226
rect 291306 4170 291374 4226
rect 291430 4170 291498 4226
rect 291554 4170 291622 4226
rect 291678 4170 291774 4226
rect 291154 4102 291774 4170
rect 291154 4046 291250 4102
rect 291306 4046 291374 4102
rect 291430 4046 291498 4102
rect 291554 4046 291622 4102
rect 291678 4046 291774 4102
rect 291154 3978 291774 4046
rect 291154 3922 291250 3978
rect 291306 3922 291374 3978
rect 291430 3922 291498 3978
rect 291554 3922 291622 3978
rect 291678 3922 291774 3978
rect 291154 -160 291774 3922
rect 291154 -216 291250 -160
rect 291306 -216 291374 -160
rect 291430 -216 291498 -160
rect 291554 -216 291622 -160
rect 291678 -216 291774 -160
rect 291154 -284 291774 -216
rect 291154 -340 291250 -284
rect 291306 -340 291374 -284
rect 291430 -340 291498 -284
rect 291554 -340 291622 -284
rect 291678 -340 291774 -284
rect 291154 -408 291774 -340
rect 291154 -464 291250 -408
rect 291306 -464 291374 -408
rect 291430 -464 291498 -408
rect 291554 -464 291622 -408
rect 291678 -464 291774 -408
rect 291154 -532 291774 -464
rect 291154 -588 291250 -532
rect 291306 -588 291374 -532
rect 291430 -588 291498 -532
rect 291554 -588 291622 -532
rect 291678 -588 291774 -532
rect 291154 -1644 291774 -588
rect 294874 28350 295494 32890
rect 294874 28294 294970 28350
rect 295026 28294 295094 28350
rect 295150 28294 295218 28350
rect 295274 28294 295342 28350
rect 295398 28294 295494 28350
rect 294874 28226 295494 28294
rect 294874 28170 294970 28226
rect 295026 28170 295094 28226
rect 295150 28170 295218 28226
rect 295274 28170 295342 28226
rect 295398 28170 295494 28226
rect 294874 28102 295494 28170
rect 294874 28046 294970 28102
rect 295026 28046 295094 28102
rect 295150 28046 295218 28102
rect 295274 28046 295342 28102
rect 295398 28046 295494 28102
rect 294874 27978 295494 28046
rect 294874 27922 294970 27978
rect 295026 27922 295094 27978
rect 295150 27922 295218 27978
rect 295274 27922 295342 27978
rect 295398 27922 295494 27978
rect 294874 10350 295494 27922
rect 294874 10294 294970 10350
rect 295026 10294 295094 10350
rect 295150 10294 295218 10350
rect 295274 10294 295342 10350
rect 295398 10294 295494 10350
rect 294874 10226 295494 10294
rect 294874 10170 294970 10226
rect 295026 10170 295094 10226
rect 295150 10170 295218 10226
rect 295274 10170 295342 10226
rect 295398 10170 295494 10226
rect 294874 10102 295494 10170
rect 294874 10046 294970 10102
rect 295026 10046 295094 10102
rect 295150 10046 295218 10102
rect 295274 10046 295342 10102
rect 295398 10046 295494 10102
rect 294874 9978 295494 10046
rect 294874 9922 294970 9978
rect 295026 9922 295094 9978
rect 295150 9922 295218 9978
rect 295274 9922 295342 9978
rect 295398 9922 295494 9978
rect 294874 -1120 295494 9922
rect 294874 -1176 294970 -1120
rect 295026 -1176 295094 -1120
rect 295150 -1176 295218 -1120
rect 295274 -1176 295342 -1120
rect 295398 -1176 295494 -1120
rect 294874 -1244 295494 -1176
rect 294874 -1300 294970 -1244
rect 295026 -1300 295094 -1244
rect 295150 -1300 295218 -1244
rect 295274 -1300 295342 -1244
rect 295398 -1300 295494 -1244
rect 294874 -1368 295494 -1300
rect 294874 -1424 294970 -1368
rect 295026 -1424 295094 -1368
rect 295150 -1424 295218 -1368
rect 295274 -1424 295342 -1368
rect 295398 -1424 295494 -1368
rect 294874 -1492 295494 -1424
rect 294874 -1548 294970 -1492
rect 295026 -1548 295094 -1492
rect 295150 -1548 295218 -1492
rect 295274 -1548 295342 -1492
rect 295398 -1548 295494 -1492
rect 294874 -1644 295494 -1548
rect 309154 22350 309774 32890
rect 309154 22294 309250 22350
rect 309306 22294 309374 22350
rect 309430 22294 309498 22350
rect 309554 22294 309622 22350
rect 309678 22294 309774 22350
rect 309154 22226 309774 22294
rect 309154 22170 309250 22226
rect 309306 22170 309374 22226
rect 309430 22170 309498 22226
rect 309554 22170 309622 22226
rect 309678 22170 309774 22226
rect 309154 22102 309774 22170
rect 309154 22046 309250 22102
rect 309306 22046 309374 22102
rect 309430 22046 309498 22102
rect 309554 22046 309622 22102
rect 309678 22046 309774 22102
rect 309154 21978 309774 22046
rect 309154 21922 309250 21978
rect 309306 21922 309374 21978
rect 309430 21922 309498 21978
rect 309554 21922 309622 21978
rect 309678 21922 309774 21978
rect 309154 4350 309774 21922
rect 309154 4294 309250 4350
rect 309306 4294 309374 4350
rect 309430 4294 309498 4350
rect 309554 4294 309622 4350
rect 309678 4294 309774 4350
rect 309154 4226 309774 4294
rect 309154 4170 309250 4226
rect 309306 4170 309374 4226
rect 309430 4170 309498 4226
rect 309554 4170 309622 4226
rect 309678 4170 309774 4226
rect 309154 4102 309774 4170
rect 309154 4046 309250 4102
rect 309306 4046 309374 4102
rect 309430 4046 309498 4102
rect 309554 4046 309622 4102
rect 309678 4046 309774 4102
rect 309154 3978 309774 4046
rect 309154 3922 309250 3978
rect 309306 3922 309374 3978
rect 309430 3922 309498 3978
rect 309554 3922 309622 3978
rect 309678 3922 309774 3978
rect 309154 -160 309774 3922
rect 309154 -216 309250 -160
rect 309306 -216 309374 -160
rect 309430 -216 309498 -160
rect 309554 -216 309622 -160
rect 309678 -216 309774 -160
rect 309154 -284 309774 -216
rect 309154 -340 309250 -284
rect 309306 -340 309374 -284
rect 309430 -340 309498 -284
rect 309554 -340 309622 -284
rect 309678 -340 309774 -284
rect 309154 -408 309774 -340
rect 309154 -464 309250 -408
rect 309306 -464 309374 -408
rect 309430 -464 309498 -408
rect 309554 -464 309622 -408
rect 309678 -464 309774 -408
rect 309154 -532 309774 -464
rect 309154 -588 309250 -532
rect 309306 -588 309374 -532
rect 309430 -588 309498 -532
rect 309554 -588 309622 -532
rect 309678 -588 309774 -532
rect 309154 -1644 309774 -588
rect 312874 28350 313494 32890
rect 312874 28294 312970 28350
rect 313026 28294 313094 28350
rect 313150 28294 313218 28350
rect 313274 28294 313342 28350
rect 313398 28294 313494 28350
rect 312874 28226 313494 28294
rect 312874 28170 312970 28226
rect 313026 28170 313094 28226
rect 313150 28170 313218 28226
rect 313274 28170 313342 28226
rect 313398 28170 313494 28226
rect 312874 28102 313494 28170
rect 312874 28046 312970 28102
rect 313026 28046 313094 28102
rect 313150 28046 313218 28102
rect 313274 28046 313342 28102
rect 313398 28046 313494 28102
rect 312874 27978 313494 28046
rect 312874 27922 312970 27978
rect 313026 27922 313094 27978
rect 313150 27922 313218 27978
rect 313274 27922 313342 27978
rect 313398 27922 313494 27978
rect 312874 10350 313494 27922
rect 312874 10294 312970 10350
rect 313026 10294 313094 10350
rect 313150 10294 313218 10350
rect 313274 10294 313342 10350
rect 313398 10294 313494 10350
rect 312874 10226 313494 10294
rect 312874 10170 312970 10226
rect 313026 10170 313094 10226
rect 313150 10170 313218 10226
rect 313274 10170 313342 10226
rect 313398 10170 313494 10226
rect 312874 10102 313494 10170
rect 312874 10046 312970 10102
rect 313026 10046 313094 10102
rect 313150 10046 313218 10102
rect 313274 10046 313342 10102
rect 313398 10046 313494 10102
rect 312874 9978 313494 10046
rect 312874 9922 312970 9978
rect 313026 9922 313094 9978
rect 313150 9922 313218 9978
rect 313274 9922 313342 9978
rect 313398 9922 313494 9978
rect 312874 -1120 313494 9922
rect 312874 -1176 312970 -1120
rect 313026 -1176 313094 -1120
rect 313150 -1176 313218 -1120
rect 313274 -1176 313342 -1120
rect 313398 -1176 313494 -1120
rect 312874 -1244 313494 -1176
rect 312874 -1300 312970 -1244
rect 313026 -1300 313094 -1244
rect 313150 -1300 313218 -1244
rect 313274 -1300 313342 -1244
rect 313398 -1300 313494 -1244
rect 312874 -1368 313494 -1300
rect 312874 -1424 312970 -1368
rect 313026 -1424 313094 -1368
rect 313150 -1424 313218 -1368
rect 313274 -1424 313342 -1368
rect 313398 -1424 313494 -1368
rect 312874 -1492 313494 -1424
rect 312874 -1548 312970 -1492
rect 313026 -1548 313094 -1492
rect 313150 -1548 313218 -1492
rect 313274 -1548 313342 -1492
rect 313398 -1548 313494 -1492
rect 312874 -1644 313494 -1548
rect 327154 22350 327774 32890
rect 327154 22294 327250 22350
rect 327306 22294 327374 22350
rect 327430 22294 327498 22350
rect 327554 22294 327622 22350
rect 327678 22294 327774 22350
rect 327154 22226 327774 22294
rect 327154 22170 327250 22226
rect 327306 22170 327374 22226
rect 327430 22170 327498 22226
rect 327554 22170 327622 22226
rect 327678 22170 327774 22226
rect 327154 22102 327774 22170
rect 327154 22046 327250 22102
rect 327306 22046 327374 22102
rect 327430 22046 327498 22102
rect 327554 22046 327622 22102
rect 327678 22046 327774 22102
rect 327154 21978 327774 22046
rect 327154 21922 327250 21978
rect 327306 21922 327374 21978
rect 327430 21922 327498 21978
rect 327554 21922 327622 21978
rect 327678 21922 327774 21978
rect 327154 4350 327774 21922
rect 327154 4294 327250 4350
rect 327306 4294 327374 4350
rect 327430 4294 327498 4350
rect 327554 4294 327622 4350
rect 327678 4294 327774 4350
rect 327154 4226 327774 4294
rect 327154 4170 327250 4226
rect 327306 4170 327374 4226
rect 327430 4170 327498 4226
rect 327554 4170 327622 4226
rect 327678 4170 327774 4226
rect 327154 4102 327774 4170
rect 327154 4046 327250 4102
rect 327306 4046 327374 4102
rect 327430 4046 327498 4102
rect 327554 4046 327622 4102
rect 327678 4046 327774 4102
rect 327154 3978 327774 4046
rect 327154 3922 327250 3978
rect 327306 3922 327374 3978
rect 327430 3922 327498 3978
rect 327554 3922 327622 3978
rect 327678 3922 327774 3978
rect 327154 -160 327774 3922
rect 327154 -216 327250 -160
rect 327306 -216 327374 -160
rect 327430 -216 327498 -160
rect 327554 -216 327622 -160
rect 327678 -216 327774 -160
rect 327154 -284 327774 -216
rect 327154 -340 327250 -284
rect 327306 -340 327374 -284
rect 327430 -340 327498 -284
rect 327554 -340 327622 -284
rect 327678 -340 327774 -284
rect 327154 -408 327774 -340
rect 327154 -464 327250 -408
rect 327306 -464 327374 -408
rect 327430 -464 327498 -408
rect 327554 -464 327622 -408
rect 327678 -464 327774 -408
rect 327154 -532 327774 -464
rect 327154 -588 327250 -532
rect 327306 -588 327374 -532
rect 327430 -588 327498 -532
rect 327554 -588 327622 -532
rect 327678 -588 327774 -532
rect 327154 -1644 327774 -588
rect 330874 28350 331494 31020
rect 330874 28294 330970 28350
rect 331026 28294 331094 28350
rect 331150 28294 331218 28350
rect 331274 28294 331342 28350
rect 331398 28294 331494 28350
rect 330874 28226 331494 28294
rect 330874 28170 330970 28226
rect 331026 28170 331094 28226
rect 331150 28170 331218 28226
rect 331274 28170 331342 28226
rect 331398 28170 331494 28226
rect 330874 28102 331494 28170
rect 330874 28046 330970 28102
rect 331026 28046 331094 28102
rect 331150 28046 331218 28102
rect 331274 28046 331342 28102
rect 331398 28046 331494 28102
rect 330874 27978 331494 28046
rect 330874 27922 330970 27978
rect 331026 27922 331094 27978
rect 331150 27922 331218 27978
rect 331274 27922 331342 27978
rect 331398 27922 331494 27978
rect 330874 10350 331494 27922
rect 330874 10294 330970 10350
rect 331026 10294 331094 10350
rect 331150 10294 331218 10350
rect 331274 10294 331342 10350
rect 331398 10294 331494 10350
rect 330874 10226 331494 10294
rect 330874 10170 330970 10226
rect 331026 10170 331094 10226
rect 331150 10170 331218 10226
rect 331274 10170 331342 10226
rect 331398 10170 331494 10226
rect 330874 10102 331494 10170
rect 330874 10046 330970 10102
rect 331026 10046 331094 10102
rect 331150 10046 331218 10102
rect 331274 10046 331342 10102
rect 331398 10046 331494 10102
rect 330874 9978 331494 10046
rect 330874 9922 330970 9978
rect 331026 9922 331094 9978
rect 331150 9922 331218 9978
rect 331274 9922 331342 9978
rect 331398 9922 331494 9978
rect 330874 -1120 331494 9922
rect 330874 -1176 330970 -1120
rect 331026 -1176 331094 -1120
rect 331150 -1176 331218 -1120
rect 331274 -1176 331342 -1120
rect 331398 -1176 331494 -1120
rect 330874 -1244 331494 -1176
rect 330874 -1300 330970 -1244
rect 331026 -1300 331094 -1244
rect 331150 -1300 331218 -1244
rect 331274 -1300 331342 -1244
rect 331398 -1300 331494 -1244
rect 330874 -1368 331494 -1300
rect 330874 -1424 330970 -1368
rect 331026 -1424 331094 -1368
rect 331150 -1424 331218 -1368
rect 331274 -1424 331342 -1368
rect 331398 -1424 331494 -1368
rect 330874 -1492 331494 -1424
rect 330874 -1548 330970 -1492
rect 331026 -1548 331094 -1492
rect 331150 -1548 331218 -1492
rect 331274 -1548 331342 -1492
rect 331398 -1548 331494 -1492
rect 330874 -1644 331494 -1548
rect 345154 22350 345774 32890
rect 345154 22294 345250 22350
rect 345306 22294 345374 22350
rect 345430 22294 345498 22350
rect 345554 22294 345622 22350
rect 345678 22294 345774 22350
rect 345154 22226 345774 22294
rect 345154 22170 345250 22226
rect 345306 22170 345374 22226
rect 345430 22170 345498 22226
rect 345554 22170 345622 22226
rect 345678 22170 345774 22226
rect 345154 22102 345774 22170
rect 345154 22046 345250 22102
rect 345306 22046 345374 22102
rect 345430 22046 345498 22102
rect 345554 22046 345622 22102
rect 345678 22046 345774 22102
rect 345154 21978 345774 22046
rect 345154 21922 345250 21978
rect 345306 21922 345374 21978
rect 345430 21922 345498 21978
rect 345554 21922 345622 21978
rect 345678 21922 345774 21978
rect 345154 4350 345774 21922
rect 345154 4294 345250 4350
rect 345306 4294 345374 4350
rect 345430 4294 345498 4350
rect 345554 4294 345622 4350
rect 345678 4294 345774 4350
rect 345154 4226 345774 4294
rect 345154 4170 345250 4226
rect 345306 4170 345374 4226
rect 345430 4170 345498 4226
rect 345554 4170 345622 4226
rect 345678 4170 345774 4226
rect 345154 4102 345774 4170
rect 345154 4046 345250 4102
rect 345306 4046 345374 4102
rect 345430 4046 345498 4102
rect 345554 4046 345622 4102
rect 345678 4046 345774 4102
rect 345154 3978 345774 4046
rect 345154 3922 345250 3978
rect 345306 3922 345374 3978
rect 345430 3922 345498 3978
rect 345554 3922 345622 3978
rect 345678 3922 345774 3978
rect 345154 -160 345774 3922
rect 345154 -216 345250 -160
rect 345306 -216 345374 -160
rect 345430 -216 345498 -160
rect 345554 -216 345622 -160
rect 345678 -216 345774 -160
rect 345154 -284 345774 -216
rect 345154 -340 345250 -284
rect 345306 -340 345374 -284
rect 345430 -340 345498 -284
rect 345554 -340 345622 -284
rect 345678 -340 345774 -284
rect 345154 -408 345774 -340
rect 345154 -464 345250 -408
rect 345306 -464 345374 -408
rect 345430 -464 345498 -408
rect 345554 -464 345622 -408
rect 345678 -464 345774 -408
rect 345154 -532 345774 -464
rect 345154 -588 345250 -532
rect 345306 -588 345374 -532
rect 345430 -588 345498 -532
rect 345554 -588 345622 -532
rect 345678 -588 345774 -532
rect 345154 -1644 345774 -588
rect 348874 28350 349494 32890
rect 348874 28294 348970 28350
rect 349026 28294 349094 28350
rect 349150 28294 349218 28350
rect 349274 28294 349342 28350
rect 349398 28294 349494 28350
rect 348874 28226 349494 28294
rect 348874 28170 348970 28226
rect 349026 28170 349094 28226
rect 349150 28170 349218 28226
rect 349274 28170 349342 28226
rect 349398 28170 349494 28226
rect 348874 28102 349494 28170
rect 348874 28046 348970 28102
rect 349026 28046 349094 28102
rect 349150 28046 349218 28102
rect 349274 28046 349342 28102
rect 349398 28046 349494 28102
rect 348874 27978 349494 28046
rect 348874 27922 348970 27978
rect 349026 27922 349094 27978
rect 349150 27922 349218 27978
rect 349274 27922 349342 27978
rect 349398 27922 349494 27978
rect 348874 10350 349494 27922
rect 348874 10294 348970 10350
rect 349026 10294 349094 10350
rect 349150 10294 349218 10350
rect 349274 10294 349342 10350
rect 349398 10294 349494 10350
rect 348874 10226 349494 10294
rect 348874 10170 348970 10226
rect 349026 10170 349094 10226
rect 349150 10170 349218 10226
rect 349274 10170 349342 10226
rect 349398 10170 349494 10226
rect 348874 10102 349494 10170
rect 348874 10046 348970 10102
rect 349026 10046 349094 10102
rect 349150 10046 349218 10102
rect 349274 10046 349342 10102
rect 349398 10046 349494 10102
rect 348874 9978 349494 10046
rect 348874 9922 348970 9978
rect 349026 9922 349094 9978
rect 349150 9922 349218 9978
rect 349274 9922 349342 9978
rect 349398 9922 349494 9978
rect 348874 -1120 349494 9922
rect 348874 -1176 348970 -1120
rect 349026 -1176 349094 -1120
rect 349150 -1176 349218 -1120
rect 349274 -1176 349342 -1120
rect 349398 -1176 349494 -1120
rect 348874 -1244 349494 -1176
rect 348874 -1300 348970 -1244
rect 349026 -1300 349094 -1244
rect 349150 -1300 349218 -1244
rect 349274 -1300 349342 -1244
rect 349398 -1300 349494 -1244
rect 348874 -1368 349494 -1300
rect 348874 -1424 348970 -1368
rect 349026 -1424 349094 -1368
rect 349150 -1424 349218 -1368
rect 349274 -1424 349342 -1368
rect 349398 -1424 349494 -1368
rect 348874 -1492 349494 -1424
rect 348874 -1548 348970 -1492
rect 349026 -1548 349094 -1492
rect 349150 -1548 349218 -1492
rect 349274 -1548 349342 -1492
rect 349398 -1548 349494 -1492
rect 348874 -1644 349494 -1548
rect 363154 22350 363774 32890
rect 363154 22294 363250 22350
rect 363306 22294 363374 22350
rect 363430 22294 363498 22350
rect 363554 22294 363622 22350
rect 363678 22294 363774 22350
rect 363154 22226 363774 22294
rect 363154 22170 363250 22226
rect 363306 22170 363374 22226
rect 363430 22170 363498 22226
rect 363554 22170 363622 22226
rect 363678 22170 363774 22226
rect 363154 22102 363774 22170
rect 363154 22046 363250 22102
rect 363306 22046 363374 22102
rect 363430 22046 363498 22102
rect 363554 22046 363622 22102
rect 363678 22046 363774 22102
rect 363154 21978 363774 22046
rect 363154 21922 363250 21978
rect 363306 21922 363374 21978
rect 363430 21922 363498 21978
rect 363554 21922 363622 21978
rect 363678 21922 363774 21978
rect 363154 4350 363774 21922
rect 363154 4294 363250 4350
rect 363306 4294 363374 4350
rect 363430 4294 363498 4350
rect 363554 4294 363622 4350
rect 363678 4294 363774 4350
rect 363154 4226 363774 4294
rect 363154 4170 363250 4226
rect 363306 4170 363374 4226
rect 363430 4170 363498 4226
rect 363554 4170 363622 4226
rect 363678 4170 363774 4226
rect 363154 4102 363774 4170
rect 363154 4046 363250 4102
rect 363306 4046 363374 4102
rect 363430 4046 363498 4102
rect 363554 4046 363622 4102
rect 363678 4046 363774 4102
rect 363154 3978 363774 4046
rect 363154 3922 363250 3978
rect 363306 3922 363374 3978
rect 363430 3922 363498 3978
rect 363554 3922 363622 3978
rect 363678 3922 363774 3978
rect 363154 -160 363774 3922
rect 363154 -216 363250 -160
rect 363306 -216 363374 -160
rect 363430 -216 363498 -160
rect 363554 -216 363622 -160
rect 363678 -216 363774 -160
rect 363154 -284 363774 -216
rect 363154 -340 363250 -284
rect 363306 -340 363374 -284
rect 363430 -340 363498 -284
rect 363554 -340 363622 -284
rect 363678 -340 363774 -284
rect 363154 -408 363774 -340
rect 363154 -464 363250 -408
rect 363306 -464 363374 -408
rect 363430 -464 363498 -408
rect 363554 -464 363622 -408
rect 363678 -464 363774 -408
rect 363154 -532 363774 -464
rect 363154 -588 363250 -532
rect 363306 -588 363374 -532
rect 363430 -588 363498 -532
rect 363554 -588 363622 -532
rect 363678 -588 363774 -532
rect 363154 -1644 363774 -588
rect 366874 28350 367494 32890
rect 366874 28294 366970 28350
rect 367026 28294 367094 28350
rect 367150 28294 367218 28350
rect 367274 28294 367342 28350
rect 367398 28294 367494 28350
rect 366874 28226 367494 28294
rect 366874 28170 366970 28226
rect 367026 28170 367094 28226
rect 367150 28170 367218 28226
rect 367274 28170 367342 28226
rect 367398 28170 367494 28226
rect 366874 28102 367494 28170
rect 366874 28046 366970 28102
rect 367026 28046 367094 28102
rect 367150 28046 367218 28102
rect 367274 28046 367342 28102
rect 367398 28046 367494 28102
rect 366874 27978 367494 28046
rect 366874 27922 366970 27978
rect 367026 27922 367094 27978
rect 367150 27922 367218 27978
rect 367274 27922 367342 27978
rect 367398 27922 367494 27978
rect 366874 10350 367494 27922
rect 366874 10294 366970 10350
rect 367026 10294 367094 10350
rect 367150 10294 367218 10350
rect 367274 10294 367342 10350
rect 367398 10294 367494 10350
rect 366874 10226 367494 10294
rect 366874 10170 366970 10226
rect 367026 10170 367094 10226
rect 367150 10170 367218 10226
rect 367274 10170 367342 10226
rect 367398 10170 367494 10226
rect 366874 10102 367494 10170
rect 366874 10046 366970 10102
rect 367026 10046 367094 10102
rect 367150 10046 367218 10102
rect 367274 10046 367342 10102
rect 367398 10046 367494 10102
rect 366874 9978 367494 10046
rect 366874 9922 366970 9978
rect 367026 9922 367094 9978
rect 367150 9922 367218 9978
rect 367274 9922 367342 9978
rect 367398 9922 367494 9978
rect 366874 -1120 367494 9922
rect 366874 -1176 366970 -1120
rect 367026 -1176 367094 -1120
rect 367150 -1176 367218 -1120
rect 367274 -1176 367342 -1120
rect 367398 -1176 367494 -1120
rect 366874 -1244 367494 -1176
rect 366874 -1300 366970 -1244
rect 367026 -1300 367094 -1244
rect 367150 -1300 367218 -1244
rect 367274 -1300 367342 -1244
rect 367398 -1300 367494 -1244
rect 366874 -1368 367494 -1300
rect 366874 -1424 366970 -1368
rect 367026 -1424 367094 -1368
rect 367150 -1424 367218 -1368
rect 367274 -1424 367342 -1368
rect 367398 -1424 367494 -1368
rect 366874 -1492 367494 -1424
rect 366874 -1548 366970 -1492
rect 367026 -1548 367094 -1492
rect 367150 -1548 367218 -1492
rect 367274 -1548 367342 -1492
rect 367398 -1548 367494 -1492
rect 366874 -1644 367494 -1548
rect 381154 22350 381774 32890
rect 381154 22294 381250 22350
rect 381306 22294 381374 22350
rect 381430 22294 381498 22350
rect 381554 22294 381622 22350
rect 381678 22294 381774 22350
rect 381154 22226 381774 22294
rect 381154 22170 381250 22226
rect 381306 22170 381374 22226
rect 381430 22170 381498 22226
rect 381554 22170 381622 22226
rect 381678 22170 381774 22226
rect 381154 22102 381774 22170
rect 381154 22046 381250 22102
rect 381306 22046 381374 22102
rect 381430 22046 381498 22102
rect 381554 22046 381622 22102
rect 381678 22046 381774 22102
rect 381154 21978 381774 22046
rect 381154 21922 381250 21978
rect 381306 21922 381374 21978
rect 381430 21922 381498 21978
rect 381554 21922 381622 21978
rect 381678 21922 381774 21978
rect 381154 4350 381774 21922
rect 381154 4294 381250 4350
rect 381306 4294 381374 4350
rect 381430 4294 381498 4350
rect 381554 4294 381622 4350
rect 381678 4294 381774 4350
rect 381154 4226 381774 4294
rect 381154 4170 381250 4226
rect 381306 4170 381374 4226
rect 381430 4170 381498 4226
rect 381554 4170 381622 4226
rect 381678 4170 381774 4226
rect 381154 4102 381774 4170
rect 381154 4046 381250 4102
rect 381306 4046 381374 4102
rect 381430 4046 381498 4102
rect 381554 4046 381622 4102
rect 381678 4046 381774 4102
rect 381154 3978 381774 4046
rect 381154 3922 381250 3978
rect 381306 3922 381374 3978
rect 381430 3922 381498 3978
rect 381554 3922 381622 3978
rect 381678 3922 381774 3978
rect 381154 -160 381774 3922
rect 381154 -216 381250 -160
rect 381306 -216 381374 -160
rect 381430 -216 381498 -160
rect 381554 -216 381622 -160
rect 381678 -216 381774 -160
rect 381154 -284 381774 -216
rect 381154 -340 381250 -284
rect 381306 -340 381374 -284
rect 381430 -340 381498 -284
rect 381554 -340 381622 -284
rect 381678 -340 381774 -284
rect 381154 -408 381774 -340
rect 381154 -464 381250 -408
rect 381306 -464 381374 -408
rect 381430 -464 381498 -408
rect 381554 -464 381622 -408
rect 381678 -464 381774 -408
rect 381154 -532 381774 -464
rect 381154 -588 381250 -532
rect 381306 -588 381374 -532
rect 381430 -588 381498 -532
rect 381554 -588 381622 -532
rect 381678 -588 381774 -532
rect 381154 -1644 381774 -588
rect 384874 28350 385494 32890
rect 384874 28294 384970 28350
rect 385026 28294 385094 28350
rect 385150 28294 385218 28350
rect 385274 28294 385342 28350
rect 385398 28294 385494 28350
rect 384874 28226 385494 28294
rect 384874 28170 384970 28226
rect 385026 28170 385094 28226
rect 385150 28170 385218 28226
rect 385274 28170 385342 28226
rect 385398 28170 385494 28226
rect 384874 28102 385494 28170
rect 384874 28046 384970 28102
rect 385026 28046 385094 28102
rect 385150 28046 385218 28102
rect 385274 28046 385342 28102
rect 385398 28046 385494 28102
rect 384874 27978 385494 28046
rect 384874 27922 384970 27978
rect 385026 27922 385094 27978
rect 385150 27922 385218 27978
rect 385274 27922 385342 27978
rect 385398 27922 385494 27978
rect 384874 10350 385494 27922
rect 384874 10294 384970 10350
rect 385026 10294 385094 10350
rect 385150 10294 385218 10350
rect 385274 10294 385342 10350
rect 385398 10294 385494 10350
rect 384874 10226 385494 10294
rect 384874 10170 384970 10226
rect 385026 10170 385094 10226
rect 385150 10170 385218 10226
rect 385274 10170 385342 10226
rect 385398 10170 385494 10226
rect 384874 10102 385494 10170
rect 384874 10046 384970 10102
rect 385026 10046 385094 10102
rect 385150 10046 385218 10102
rect 385274 10046 385342 10102
rect 385398 10046 385494 10102
rect 384874 9978 385494 10046
rect 384874 9922 384970 9978
rect 385026 9922 385094 9978
rect 385150 9922 385218 9978
rect 385274 9922 385342 9978
rect 385398 9922 385494 9978
rect 384874 -1120 385494 9922
rect 384874 -1176 384970 -1120
rect 385026 -1176 385094 -1120
rect 385150 -1176 385218 -1120
rect 385274 -1176 385342 -1120
rect 385398 -1176 385494 -1120
rect 384874 -1244 385494 -1176
rect 384874 -1300 384970 -1244
rect 385026 -1300 385094 -1244
rect 385150 -1300 385218 -1244
rect 385274 -1300 385342 -1244
rect 385398 -1300 385494 -1244
rect 384874 -1368 385494 -1300
rect 384874 -1424 384970 -1368
rect 385026 -1424 385094 -1368
rect 385150 -1424 385218 -1368
rect 385274 -1424 385342 -1368
rect 385398 -1424 385494 -1368
rect 384874 -1492 385494 -1424
rect 384874 -1548 384970 -1492
rect 385026 -1548 385094 -1492
rect 385150 -1548 385218 -1492
rect 385274 -1548 385342 -1492
rect 385398 -1548 385494 -1492
rect 384874 -1644 385494 -1548
rect 399154 22350 399774 32890
rect 399154 22294 399250 22350
rect 399306 22294 399374 22350
rect 399430 22294 399498 22350
rect 399554 22294 399622 22350
rect 399678 22294 399774 22350
rect 399154 22226 399774 22294
rect 399154 22170 399250 22226
rect 399306 22170 399374 22226
rect 399430 22170 399498 22226
rect 399554 22170 399622 22226
rect 399678 22170 399774 22226
rect 399154 22102 399774 22170
rect 399154 22046 399250 22102
rect 399306 22046 399374 22102
rect 399430 22046 399498 22102
rect 399554 22046 399622 22102
rect 399678 22046 399774 22102
rect 399154 21978 399774 22046
rect 399154 21922 399250 21978
rect 399306 21922 399374 21978
rect 399430 21922 399498 21978
rect 399554 21922 399622 21978
rect 399678 21922 399774 21978
rect 399154 4350 399774 21922
rect 399154 4294 399250 4350
rect 399306 4294 399374 4350
rect 399430 4294 399498 4350
rect 399554 4294 399622 4350
rect 399678 4294 399774 4350
rect 399154 4226 399774 4294
rect 399154 4170 399250 4226
rect 399306 4170 399374 4226
rect 399430 4170 399498 4226
rect 399554 4170 399622 4226
rect 399678 4170 399774 4226
rect 399154 4102 399774 4170
rect 399154 4046 399250 4102
rect 399306 4046 399374 4102
rect 399430 4046 399498 4102
rect 399554 4046 399622 4102
rect 399678 4046 399774 4102
rect 399154 3978 399774 4046
rect 399154 3922 399250 3978
rect 399306 3922 399374 3978
rect 399430 3922 399498 3978
rect 399554 3922 399622 3978
rect 399678 3922 399774 3978
rect 399154 -160 399774 3922
rect 399154 -216 399250 -160
rect 399306 -216 399374 -160
rect 399430 -216 399498 -160
rect 399554 -216 399622 -160
rect 399678 -216 399774 -160
rect 399154 -284 399774 -216
rect 399154 -340 399250 -284
rect 399306 -340 399374 -284
rect 399430 -340 399498 -284
rect 399554 -340 399622 -284
rect 399678 -340 399774 -284
rect 399154 -408 399774 -340
rect 399154 -464 399250 -408
rect 399306 -464 399374 -408
rect 399430 -464 399498 -408
rect 399554 -464 399622 -408
rect 399678 -464 399774 -408
rect 399154 -532 399774 -464
rect 399154 -588 399250 -532
rect 399306 -588 399374 -532
rect 399430 -588 399498 -532
rect 399554 -588 399622 -532
rect 399678 -588 399774 -532
rect 399154 -1644 399774 -588
rect 402874 28350 403494 32890
rect 402874 28294 402970 28350
rect 403026 28294 403094 28350
rect 403150 28294 403218 28350
rect 403274 28294 403342 28350
rect 403398 28294 403494 28350
rect 402874 28226 403494 28294
rect 402874 28170 402970 28226
rect 403026 28170 403094 28226
rect 403150 28170 403218 28226
rect 403274 28170 403342 28226
rect 403398 28170 403494 28226
rect 402874 28102 403494 28170
rect 402874 28046 402970 28102
rect 403026 28046 403094 28102
rect 403150 28046 403218 28102
rect 403274 28046 403342 28102
rect 403398 28046 403494 28102
rect 402874 27978 403494 28046
rect 402874 27922 402970 27978
rect 403026 27922 403094 27978
rect 403150 27922 403218 27978
rect 403274 27922 403342 27978
rect 403398 27922 403494 27978
rect 402874 10350 403494 27922
rect 402874 10294 402970 10350
rect 403026 10294 403094 10350
rect 403150 10294 403218 10350
rect 403274 10294 403342 10350
rect 403398 10294 403494 10350
rect 402874 10226 403494 10294
rect 402874 10170 402970 10226
rect 403026 10170 403094 10226
rect 403150 10170 403218 10226
rect 403274 10170 403342 10226
rect 403398 10170 403494 10226
rect 402874 10102 403494 10170
rect 402874 10046 402970 10102
rect 403026 10046 403094 10102
rect 403150 10046 403218 10102
rect 403274 10046 403342 10102
rect 403398 10046 403494 10102
rect 402874 9978 403494 10046
rect 402874 9922 402970 9978
rect 403026 9922 403094 9978
rect 403150 9922 403218 9978
rect 403274 9922 403342 9978
rect 403398 9922 403494 9978
rect 402874 -1120 403494 9922
rect 402874 -1176 402970 -1120
rect 403026 -1176 403094 -1120
rect 403150 -1176 403218 -1120
rect 403274 -1176 403342 -1120
rect 403398 -1176 403494 -1120
rect 402874 -1244 403494 -1176
rect 402874 -1300 402970 -1244
rect 403026 -1300 403094 -1244
rect 403150 -1300 403218 -1244
rect 403274 -1300 403342 -1244
rect 403398 -1300 403494 -1244
rect 402874 -1368 403494 -1300
rect 402874 -1424 402970 -1368
rect 403026 -1424 403094 -1368
rect 403150 -1424 403218 -1368
rect 403274 -1424 403342 -1368
rect 403398 -1424 403494 -1368
rect 402874 -1492 403494 -1424
rect 402874 -1548 402970 -1492
rect 403026 -1548 403094 -1492
rect 403150 -1548 403218 -1492
rect 403274 -1548 403342 -1492
rect 403398 -1548 403494 -1492
rect 402874 -1644 403494 -1548
rect 417154 22350 417774 32890
rect 417154 22294 417250 22350
rect 417306 22294 417374 22350
rect 417430 22294 417498 22350
rect 417554 22294 417622 22350
rect 417678 22294 417774 22350
rect 417154 22226 417774 22294
rect 417154 22170 417250 22226
rect 417306 22170 417374 22226
rect 417430 22170 417498 22226
rect 417554 22170 417622 22226
rect 417678 22170 417774 22226
rect 417154 22102 417774 22170
rect 417154 22046 417250 22102
rect 417306 22046 417374 22102
rect 417430 22046 417498 22102
rect 417554 22046 417622 22102
rect 417678 22046 417774 22102
rect 417154 21978 417774 22046
rect 417154 21922 417250 21978
rect 417306 21922 417374 21978
rect 417430 21922 417498 21978
rect 417554 21922 417622 21978
rect 417678 21922 417774 21978
rect 417154 4350 417774 21922
rect 417154 4294 417250 4350
rect 417306 4294 417374 4350
rect 417430 4294 417498 4350
rect 417554 4294 417622 4350
rect 417678 4294 417774 4350
rect 417154 4226 417774 4294
rect 417154 4170 417250 4226
rect 417306 4170 417374 4226
rect 417430 4170 417498 4226
rect 417554 4170 417622 4226
rect 417678 4170 417774 4226
rect 417154 4102 417774 4170
rect 417154 4046 417250 4102
rect 417306 4046 417374 4102
rect 417430 4046 417498 4102
rect 417554 4046 417622 4102
rect 417678 4046 417774 4102
rect 417154 3978 417774 4046
rect 417154 3922 417250 3978
rect 417306 3922 417374 3978
rect 417430 3922 417498 3978
rect 417554 3922 417622 3978
rect 417678 3922 417774 3978
rect 417154 -160 417774 3922
rect 417154 -216 417250 -160
rect 417306 -216 417374 -160
rect 417430 -216 417498 -160
rect 417554 -216 417622 -160
rect 417678 -216 417774 -160
rect 417154 -284 417774 -216
rect 417154 -340 417250 -284
rect 417306 -340 417374 -284
rect 417430 -340 417498 -284
rect 417554 -340 417622 -284
rect 417678 -340 417774 -284
rect 417154 -408 417774 -340
rect 417154 -464 417250 -408
rect 417306 -464 417374 -408
rect 417430 -464 417498 -408
rect 417554 -464 417622 -408
rect 417678 -464 417774 -408
rect 417154 -532 417774 -464
rect 417154 -588 417250 -532
rect 417306 -588 417374 -532
rect 417430 -588 417498 -532
rect 417554 -588 417622 -532
rect 417678 -588 417774 -532
rect 417154 -1644 417774 -588
rect 420874 28350 421494 32890
rect 420874 28294 420970 28350
rect 421026 28294 421094 28350
rect 421150 28294 421218 28350
rect 421274 28294 421342 28350
rect 421398 28294 421494 28350
rect 420874 28226 421494 28294
rect 420874 28170 420970 28226
rect 421026 28170 421094 28226
rect 421150 28170 421218 28226
rect 421274 28170 421342 28226
rect 421398 28170 421494 28226
rect 420874 28102 421494 28170
rect 420874 28046 420970 28102
rect 421026 28046 421094 28102
rect 421150 28046 421218 28102
rect 421274 28046 421342 28102
rect 421398 28046 421494 28102
rect 420874 27978 421494 28046
rect 420874 27922 420970 27978
rect 421026 27922 421094 27978
rect 421150 27922 421218 27978
rect 421274 27922 421342 27978
rect 421398 27922 421494 27978
rect 420874 10350 421494 27922
rect 420874 10294 420970 10350
rect 421026 10294 421094 10350
rect 421150 10294 421218 10350
rect 421274 10294 421342 10350
rect 421398 10294 421494 10350
rect 420874 10226 421494 10294
rect 420874 10170 420970 10226
rect 421026 10170 421094 10226
rect 421150 10170 421218 10226
rect 421274 10170 421342 10226
rect 421398 10170 421494 10226
rect 420874 10102 421494 10170
rect 420874 10046 420970 10102
rect 421026 10046 421094 10102
rect 421150 10046 421218 10102
rect 421274 10046 421342 10102
rect 421398 10046 421494 10102
rect 420874 9978 421494 10046
rect 420874 9922 420970 9978
rect 421026 9922 421094 9978
rect 421150 9922 421218 9978
rect 421274 9922 421342 9978
rect 421398 9922 421494 9978
rect 420874 -1120 421494 9922
rect 420874 -1176 420970 -1120
rect 421026 -1176 421094 -1120
rect 421150 -1176 421218 -1120
rect 421274 -1176 421342 -1120
rect 421398 -1176 421494 -1120
rect 420874 -1244 421494 -1176
rect 420874 -1300 420970 -1244
rect 421026 -1300 421094 -1244
rect 421150 -1300 421218 -1244
rect 421274 -1300 421342 -1244
rect 421398 -1300 421494 -1244
rect 420874 -1368 421494 -1300
rect 420874 -1424 420970 -1368
rect 421026 -1424 421094 -1368
rect 421150 -1424 421218 -1368
rect 421274 -1424 421342 -1368
rect 421398 -1424 421494 -1368
rect 420874 -1492 421494 -1424
rect 420874 -1548 420970 -1492
rect 421026 -1548 421094 -1492
rect 421150 -1548 421218 -1492
rect 421274 -1548 421342 -1492
rect 421398 -1548 421494 -1492
rect 420874 -1644 421494 -1548
rect 435154 22350 435774 32890
rect 435154 22294 435250 22350
rect 435306 22294 435374 22350
rect 435430 22294 435498 22350
rect 435554 22294 435622 22350
rect 435678 22294 435774 22350
rect 435154 22226 435774 22294
rect 435154 22170 435250 22226
rect 435306 22170 435374 22226
rect 435430 22170 435498 22226
rect 435554 22170 435622 22226
rect 435678 22170 435774 22226
rect 435154 22102 435774 22170
rect 435154 22046 435250 22102
rect 435306 22046 435374 22102
rect 435430 22046 435498 22102
rect 435554 22046 435622 22102
rect 435678 22046 435774 22102
rect 435154 21978 435774 22046
rect 435154 21922 435250 21978
rect 435306 21922 435374 21978
rect 435430 21922 435498 21978
rect 435554 21922 435622 21978
rect 435678 21922 435774 21978
rect 435154 4350 435774 21922
rect 435154 4294 435250 4350
rect 435306 4294 435374 4350
rect 435430 4294 435498 4350
rect 435554 4294 435622 4350
rect 435678 4294 435774 4350
rect 435154 4226 435774 4294
rect 435154 4170 435250 4226
rect 435306 4170 435374 4226
rect 435430 4170 435498 4226
rect 435554 4170 435622 4226
rect 435678 4170 435774 4226
rect 435154 4102 435774 4170
rect 435154 4046 435250 4102
rect 435306 4046 435374 4102
rect 435430 4046 435498 4102
rect 435554 4046 435622 4102
rect 435678 4046 435774 4102
rect 435154 3978 435774 4046
rect 435154 3922 435250 3978
rect 435306 3922 435374 3978
rect 435430 3922 435498 3978
rect 435554 3922 435622 3978
rect 435678 3922 435774 3978
rect 435154 -160 435774 3922
rect 435154 -216 435250 -160
rect 435306 -216 435374 -160
rect 435430 -216 435498 -160
rect 435554 -216 435622 -160
rect 435678 -216 435774 -160
rect 435154 -284 435774 -216
rect 435154 -340 435250 -284
rect 435306 -340 435374 -284
rect 435430 -340 435498 -284
rect 435554 -340 435622 -284
rect 435678 -340 435774 -284
rect 435154 -408 435774 -340
rect 435154 -464 435250 -408
rect 435306 -464 435374 -408
rect 435430 -464 435498 -408
rect 435554 -464 435622 -408
rect 435678 -464 435774 -408
rect 435154 -532 435774 -464
rect 435154 -588 435250 -532
rect 435306 -588 435374 -532
rect 435430 -588 435498 -532
rect 435554 -588 435622 -532
rect 435678 -588 435774 -532
rect 435154 -1644 435774 -588
rect 438874 28350 439494 32890
rect 438874 28294 438970 28350
rect 439026 28294 439094 28350
rect 439150 28294 439218 28350
rect 439274 28294 439342 28350
rect 439398 28294 439494 28350
rect 438874 28226 439494 28294
rect 438874 28170 438970 28226
rect 439026 28170 439094 28226
rect 439150 28170 439218 28226
rect 439274 28170 439342 28226
rect 439398 28170 439494 28226
rect 438874 28102 439494 28170
rect 438874 28046 438970 28102
rect 439026 28046 439094 28102
rect 439150 28046 439218 28102
rect 439274 28046 439342 28102
rect 439398 28046 439494 28102
rect 438874 27978 439494 28046
rect 438874 27922 438970 27978
rect 439026 27922 439094 27978
rect 439150 27922 439218 27978
rect 439274 27922 439342 27978
rect 439398 27922 439494 27978
rect 438874 10350 439494 27922
rect 438874 10294 438970 10350
rect 439026 10294 439094 10350
rect 439150 10294 439218 10350
rect 439274 10294 439342 10350
rect 439398 10294 439494 10350
rect 438874 10226 439494 10294
rect 438874 10170 438970 10226
rect 439026 10170 439094 10226
rect 439150 10170 439218 10226
rect 439274 10170 439342 10226
rect 439398 10170 439494 10226
rect 438874 10102 439494 10170
rect 438874 10046 438970 10102
rect 439026 10046 439094 10102
rect 439150 10046 439218 10102
rect 439274 10046 439342 10102
rect 439398 10046 439494 10102
rect 438874 9978 439494 10046
rect 438874 9922 438970 9978
rect 439026 9922 439094 9978
rect 439150 9922 439218 9978
rect 439274 9922 439342 9978
rect 439398 9922 439494 9978
rect 438874 -1120 439494 9922
rect 438874 -1176 438970 -1120
rect 439026 -1176 439094 -1120
rect 439150 -1176 439218 -1120
rect 439274 -1176 439342 -1120
rect 439398 -1176 439494 -1120
rect 438874 -1244 439494 -1176
rect 438874 -1300 438970 -1244
rect 439026 -1300 439094 -1244
rect 439150 -1300 439218 -1244
rect 439274 -1300 439342 -1244
rect 439398 -1300 439494 -1244
rect 438874 -1368 439494 -1300
rect 438874 -1424 438970 -1368
rect 439026 -1424 439094 -1368
rect 439150 -1424 439218 -1368
rect 439274 -1424 439342 -1368
rect 439398 -1424 439494 -1368
rect 438874 -1492 439494 -1424
rect 438874 -1548 438970 -1492
rect 439026 -1548 439094 -1492
rect 439150 -1548 439218 -1492
rect 439274 -1548 439342 -1492
rect 439398 -1548 439494 -1492
rect 438874 -1644 439494 -1548
rect 453154 22350 453774 31020
rect 453154 22294 453250 22350
rect 453306 22294 453374 22350
rect 453430 22294 453498 22350
rect 453554 22294 453622 22350
rect 453678 22294 453774 22350
rect 453154 22226 453774 22294
rect 453154 22170 453250 22226
rect 453306 22170 453374 22226
rect 453430 22170 453498 22226
rect 453554 22170 453622 22226
rect 453678 22170 453774 22226
rect 453154 22102 453774 22170
rect 453154 22046 453250 22102
rect 453306 22046 453374 22102
rect 453430 22046 453498 22102
rect 453554 22046 453622 22102
rect 453678 22046 453774 22102
rect 453154 21978 453774 22046
rect 453154 21922 453250 21978
rect 453306 21922 453374 21978
rect 453430 21922 453498 21978
rect 453554 21922 453622 21978
rect 453678 21922 453774 21978
rect 453154 4350 453774 21922
rect 453154 4294 453250 4350
rect 453306 4294 453374 4350
rect 453430 4294 453498 4350
rect 453554 4294 453622 4350
rect 453678 4294 453774 4350
rect 453154 4226 453774 4294
rect 453154 4170 453250 4226
rect 453306 4170 453374 4226
rect 453430 4170 453498 4226
rect 453554 4170 453622 4226
rect 453678 4170 453774 4226
rect 453154 4102 453774 4170
rect 453154 4046 453250 4102
rect 453306 4046 453374 4102
rect 453430 4046 453498 4102
rect 453554 4046 453622 4102
rect 453678 4046 453774 4102
rect 453154 3978 453774 4046
rect 453154 3922 453250 3978
rect 453306 3922 453374 3978
rect 453430 3922 453498 3978
rect 453554 3922 453622 3978
rect 453678 3922 453774 3978
rect 453154 -160 453774 3922
rect 453154 -216 453250 -160
rect 453306 -216 453374 -160
rect 453430 -216 453498 -160
rect 453554 -216 453622 -160
rect 453678 -216 453774 -160
rect 453154 -284 453774 -216
rect 453154 -340 453250 -284
rect 453306 -340 453374 -284
rect 453430 -340 453498 -284
rect 453554 -340 453622 -284
rect 453678 -340 453774 -284
rect 453154 -408 453774 -340
rect 453154 -464 453250 -408
rect 453306 -464 453374 -408
rect 453430 -464 453498 -408
rect 453554 -464 453622 -408
rect 453678 -464 453774 -408
rect 453154 -532 453774 -464
rect 453154 -588 453250 -532
rect 453306 -588 453374 -532
rect 453430 -588 453498 -532
rect 453554 -588 453622 -532
rect 453678 -588 453774 -532
rect 453154 -1644 453774 -588
rect 456874 28350 457494 32890
rect 456874 28294 456970 28350
rect 457026 28294 457094 28350
rect 457150 28294 457218 28350
rect 457274 28294 457342 28350
rect 457398 28294 457494 28350
rect 456874 28226 457494 28294
rect 456874 28170 456970 28226
rect 457026 28170 457094 28226
rect 457150 28170 457218 28226
rect 457274 28170 457342 28226
rect 457398 28170 457494 28226
rect 456874 28102 457494 28170
rect 456874 28046 456970 28102
rect 457026 28046 457094 28102
rect 457150 28046 457218 28102
rect 457274 28046 457342 28102
rect 457398 28046 457494 28102
rect 456874 27978 457494 28046
rect 456874 27922 456970 27978
rect 457026 27922 457094 27978
rect 457150 27922 457218 27978
rect 457274 27922 457342 27978
rect 457398 27922 457494 27978
rect 456874 10350 457494 27922
rect 456874 10294 456970 10350
rect 457026 10294 457094 10350
rect 457150 10294 457218 10350
rect 457274 10294 457342 10350
rect 457398 10294 457494 10350
rect 456874 10226 457494 10294
rect 456874 10170 456970 10226
rect 457026 10170 457094 10226
rect 457150 10170 457218 10226
rect 457274 10170 457342 10226
rect 457398 10170 457494 10226
rect 456874 10102 457494 10170
rect 456874 10046 456970 10102
rect 457026 10046 457094 10102
rect 457150 10046 457218 10102
rect 457274 10046 457342 10102
rect 457398 10046 457494 10102
rect 456874 9978 457494 10046
rect 456874 9922 456970 9978
rect 457026 9922 457094 9978
rect 457150 9922 457218 9978
rect 457274 9922 457342 9978
rect 457398 9922 457494 9978
rect 456874 -1120 457494 9922
rect 456874 -1176 456970 -1120
rect 457026 -1176 457094 -1120
rect 457150 -1176 457218 -1120
rect 457274 -1176 457342 -1120
rect 457398 -1176 457494 -1120
rect 456874 -1244 457494 -1176
rect 456874 -1300 456970 -1244
rect 457026 -1300 457094 -1244
rect 457150 -1300 457218 -1244
rect 457274 -1300 457342 -1244
rect 457398 -1300 457494 -1244
rect 456874 -1368 457494 -1300
rect 456874 -1424 456970 -1368
rect 457026 -1424 457094 -1368
rect 457150 -1424 457218 -1368
rect 457274 -1424 457342 -1368
rect 457398 -1424 457494 -1368
rect 456874 -1492 457494 -1424
rect 456874 -1548 456970 -1492
rect 457026 -1548 457094 -1492
rect 457150 -1548 457218 -1492
rect 457274 -1548 457342 -1492
rect 457398 -1548 457494 -1492
rect 456874 -1644 457494 -1548
rect 471154 22350 471774 32890
rect 471154 22294 471250 22350
rect 471306 22294 471374 22350
rect 471430 22294 471498 22350
rect 471554 22294 471622 22350
rect 471678 22294 471774 22350
rect 471154 22226 471774 22294
rect 471154 22170 471250 22226
rect 471306 22170 471374 22226
rect 471430 22170 471498 22226
rect 471554 22170 471622 22226
rect 471678 22170 471774 22226
rect 471154 22102 471774 22170
rect 471154 22046 471250 22102
rect 471306 22046 471374 22102
rect 471430 22046 471498 22102
rect 471554 22046 471622 22102
rect 471678 22046 471774 22102
rect 471154 21978 471774 22046
rect 471154 21922 471250 21978
rect 471306 21922 471374 21978
rect 471430 21922 471498 21978
rect 471554 21922 471622 21978
rect 471678 21922 471774 21978
rect 471154 4350 471774 21922
rect 471154 4294 471250 4350
rect 471306 4294 471374 4350
rect 471430 4294 471498 4350
rect 471554 4294 471622 4350
rect 471678 4294 471774 4350
rect 471154 4226 471774 4294
rect 471154 4170 471250 4226
rect 471306 4170 471374 4226
rect 471430 4170 471498 4226
rect 471554 4170 471622 4226
rect 471678 4170 471774 4226
rect 471154 4102 471774 4170
rect 471154 4046 471250 4102
rect 471306 4046 471374 4102
rect 471430 4046 471498 4102
rect 471554 4046 471622 4102
rect 471678 4046 471774 4102
rect 471154 3978 471774 4046
rect 471154 3922 471250 3978
rect 471306 3922 471374 3978
rect 471430 3922 471498 3978
rect 471554 3922 471622 3978
rect 471678 3922 471774 3978
rect 471154 -160 471774 3922
rect 471154 -216 471250 -160
rect 471306 -216 471374 -160
rect 471430 -216 471498 -160
rect 471554 -216 471622 -160
rect 471678 -216 471774 -160
rect 471154 -284 471774 -216
rect 471154 -340 471250 -284
rect 471306 -340 471374 -284
rect 471430 -340 471498 -284
rect 471554 -340 471622 -284
rect 471678 -340 471774 -284
rect 471154 -408 471774 -340
rect 471154 -464 471250 -408
rect 471306 -464 471374 -408
rect 471430 -464 471498 -408
rect 471554 -464 471622 -408
rect 471678 -464 471774 -408
rect 471154 -532 471774 -464
rect 471154 -588 471250 -532
rect 471306 -588 471374 -532
rect 471430 -588 471498 -532
rect 471554 -588 471622 -532
rect 471678 -588 471774 -532
rect 471154 -1644 471774 -588
rect 474874 28350 475494 32890
rect 474874 28294 474970 28350
rect 475026 28294 475094 28350
rect 475150 28294 475218 28350
rect 475274 28294 475342 28350
rect 475398 28294 475494 28350
rect 474874 28226 475494 28294
rect 474874 28170 474970 28226
rect 475026 28170 475094 28226
rect 475150 28170 475218 28226
rect 475274 28170 475342 28226
rect 475398 28170 475494 28226
rect 474874 28102 475494 28170
rect 474874 28046 474970 28102
rect 475026 28046 475094 28102
rect 475150 28046 475218 28102
rect 475274 28046 475342 28102
rect 475398 28046 475494 28102
rect 474874 27978 475494 28046
rect 474874 27922 474970 27978
rect 475026 27922 475094 27978
rect 475150 27922 475218 27978
rect 475274 27922 475342 27978
rect 475398 27922 475494 27978
rect 474874 10350 475494 27922
rect 474874 10294 474970 10350
rect 475026 10294 475094 10350
rect 475150 10294 475218 10350
rect 475274 10294 475342 10350
rect 475398 10294 475494 10350
rect 474874 10226 475494 10294
rect 474874 10170 474970 10226
rect 475026 10170 475094 10226
rect 475150 10170 475218 10226
rect 475274 10170 475342 10226
rect 475398 10170 475494 10226
rect 474874 10102 475494 10170
rect 474874 10046 474970 10102
rect 475026 10046 475094 10102
rect 475150 10046 475218 10102
rect 475274 10046 475342 10102
rect 475398 10046 475494 10102
rect 474874 9978 475494 10046
rect 474874 9922 474970 9978
rect 475026 9922 475094 9978
rect 475150 9922 475218 9978
rect 475274 9922 475342 9978
rect 475398 9922 475494 9978
rect 474874 -1120 475494 9922
rect 474874 -1176 474970 -1120
rect 475026 -1176 475094 -1120
rect 475150 -1176 475218 -1120
rect 475274 -1176 475342 -1120
rect 475398 -1176 475494 -1120
rect 474874 -1244 475494 -1176
rect 474874 -1300 474970 -1244
rect 475026 -1300 475094 -1244
rect 475150 -1300 475218 -1244
rect 475274 -1300 475342 -1244
rect 475398 -1300 475494 -1244
rect 474874 -1368 475494 -1300
rect 474874 -1424 474970 -1368
rect 475026 -1424 475094 -1368
rect 475150 -1424 475218 -1368
rect 475274 -1424 475342 -1368
rect 475398 -1424 475494 -1368
rect 474874 -1492 475494 -1424
rect 474874 -1548 474970 -1492
rect 475026 -1548 475094 -1492
rect 475150 -1548 475218 -1492
rect 475274 -1548 475342 -1492
rect 475398 -1548 475494 -1492
rect 474874 -1644 475494 -1548
rect 489154 22350 489774 32890
rect 489154 22294 489250 22350
rect 489306 22294 489374 22350
rect 489430 22294 489498 22350
rect 489554 22294 489622 22350
rect 489678 22294 489774 22350
rect 489154 22226 489774 22294
rect 489154 22170 489250 22226
rect 489306 22170 489374 22226
rect 489430 22170 489498 22226
rect 489554 22170 489622 22226
rect 489678 22170 489774 22226
rect 489154 22102 489774 22170
rect 489154 22046 489250 22102
rect 489306 22046 489374 22102
rect 489430 22046 489498 22102
rect 489554 22046 489622 22102
rect 489678 22046 489774 22102
rect 489154 21978 489774 22046
rect 489154 21922 489250 21978
rect 489306 21922 489374 21978
rect 489430 21922 489498 21978
rect 489554 21922 489622 21978
rect 489678 21922 489774 21978
rect 489154 4350 489774 21922
rect 489154 4294 489250 4350
rect 489306 4294 489374 4350
rect 489430 4294 489498 4350
rect 489554 4294 489622 4350
rect 489678 4294 489774 4350
rect 489154 4226 489774 4294
rect 489154 4170 489250 4226
rect 489306 4170 489374 4226
rect 489430 4170 489498 4226
rect 489554 4170 489622 4226
rect 489678 4170 489774 4226
rect 489154 4102 489774 4170
rect 489154 4046 489250 4102
rect 489306 4046 489374 4102
rect 489430 4046 489498 4102
rect 489554 4046 489622 4102
rect 489678 4046 489774 4102
rect 489154 3978 489774 4046
rect 489154 3922 489250 3978
rect 489306 3922 489374 3978
rect 489430 3922 489498 3978
rect 489554 3922 489622 3978
rect 489678 3922 489774 3978
rect 489154 -160 489774 3922
rect 489154 -216 489250 -160
rect 489306 -216 489374 -160
rect 489430 -216 489498 -160
rect 489554 -216 489622 -160
rect 489678 -216 489774 -160
rect 489154 -284 489774 -216
rect 489154 -340 489250 -284
rect 489306 -340 489374 -284
rect 489430 -340 489498 -284
rect 489554 -340 489622 -284
rect 489678 -340 489774 -284
rect 489154 -408 489774 -340
rect 489154 -464 489250 -408
rect 489306 -464 489374 -408
rect 489430 -464 489498 -408
rect 489554 -464 489622 -408
rect 489678 -464 489774 -408
rect 489154 -532 489774 -464
rect 489154 -588 489250 -532
rect 489306 -588 489374 -532
rect 489430 -588 489498 -532
rect 489554 -588 489622 -532
rect 489678 -588 489774 -532
rect 489154 -1644 489774 -588
rect 492874 28350 493494 32890
rect 492874 28294 492970 28350
rect 493026 28294 493094 28350
rect 493150 28294 493218 28350
rect 493274 28294 493342 28350
rect 493398 28294 493494 28350
rect 492874 28226 493494 28294
rect 492874 28170 492970 28226
rect 493026 28170 493094 28226
rect 493150 28170 493218 28226
rect 493274 28170 493342 28226
rect 493398 28170 493494 28226
rect 492874 28102 493494 28170
rect 492874 28046 492970 28102
rect 493026 28046 493094 28102
rect 493150 28046 493218 28102
rect 493274 28046 493342 28102
rect 493398 28046 493494 28102
rect 492874 27978 493494 28046
rect 492874 27922 492970 27978
rect 493026 27922 493094 27978
rect 493150 27922 493218 27978
rect 493274 27922 493342 27978
rect 493398 27922 493494 27978
rect 492874 10350 493494 27922
rect 492874 10294 492970 10350
rect 493026 10294 493094 10350
rect 493150 10294 493218 10350
rect 493274 10294 493342 10350
rect 493398 10294 493494 10350
rect 492874 10226 493494 10294
rect 492874 10170 492970 10226
rect 493026 10170 493094 10226
rect 493150 10170 493218 10226
rect 493274 10170 493342 10226
rect 493398 10170 493494 10226
rect 492874 10102 493494 10170
rect 492874 10046 492970 10102
rect 493026 10046 493094 10102
rect 493150 10046 493218 10102
rect 493274 10046 493342 10102
rect 493398 10046 493494 10102
rect 492874 9978 493494 10046
rect 492874 9922 492970 9978
rect 493026 9922 493094 9978
rect 493150 9922 493218 9978
rect 493274 9922 493342 9978
rect 493398 9922 493494 9978
rect 492874 -1120 493494 9922
rect 492874 -1176 492970 -1120
rect 493026 -1176 493094 -1120
rect 493150 -1176 493218 -1120
rect 493274 -1176 493342 -1120
rect 493398 -1176 493494 -1120
rect 492874 -1244 493494 -1176
rect 492874 -1300 492970 -1244
rect 493026 -1300 493094 -1244
rect 493150 -1300 493218 -1244
rect 493274 -1300 493342 -1244
rect 493398 -1300 493494 -1244
rect 492874 -1368 493494 -1300
rect 492874 -1424 492970 -1368
rect 493026 -1424 493094 -1368
rect 493150 -1424 493218 -1368
rect 493274 -1424 493342 -1368
rect 493398 -1424 493494 -1368
rect 492874 -1492 493494 -1424
rect 492874 -1548 492970 -1492
rect 493026 -1548 493094 -1492
rect 493150 -1548 493218 -1492
rect 493274 -1548 493342 -1492
rect 493398 -1548 493494 -1492
rect 492874 -1644 493494 -1548
rect 507154 22350 507774 32890
rect 507154 22294 507250 22350
rect 507306 22294 507374 22350
rect 507430 22294 507498 22350
rect 507554 22294 507622 22350
rect 507678 22294 507774 22350
rect 507154 22226 507774 22294
rect 507154 22170 507250 22226
rect 507306 22170 507374 22226
rect 507430 22170 507498 22226
rect 507554 22170 507622 22226
rect 507678 22170 507774 22226
rect 507154 22102 507774 22170
rect 507154 22046 507250 22102
rect 507306 22046 507374 22102
rect 507430 22046 507498 22102
rect 507554 22046 507622 22102
rect 507678 22046 507774 22102
rect 507154 21978 507774 22046
rect 507154 21922 507250 21978
rect 507306 21922 507374 21978
rect 507430 21922 507498 21978
rect 507554 21922 507622 21978
rect 507678 21922 507774 21978
rect 507154 4350 507774 21922
rect 507154 4294 507250 4350
rect 507306 4294 507374 4350
rect 507430 4294 507498 4350
rect 507554 4294 507622 4350
rect 507678 4294 507774 4350
rect 507154 4226 507774 4294
rect 507154 4170 507250 4226
rect 507306 4170 507374 4226
rect 507430 4170 507498 4226
rect 507554 4170 507622 4226
rect 507678 4170 507774 4226
rect 507154 4102 507774 4170
rect 507154 4046 507250 4102
rect 507306 4046 507374 4102
rect 507430 4046 507498 4102
rect 507554 4046 507622 4102
rect 507678 4046 507774 4102
rect 507154 3978 507774 4046
rect 507154 3922 507250 3978
rect 507306 3922 507374 3978
rect 507430 3922 507498 3978
rect 507554 3922 507622 3978
rect 507678 3922 507774 3978
rect 507154 -160 507774 3922
rect 507154 -216 507250 -160
rect 507306 -216 507374 -160
rect 507430 -216 507498 -160
rect 507554 -216 507622 -160
rect 507678 -216 507774 -160
rect 507154 -284 507774 -216
rect 507154 -340 507250 -284
rect 507306 -340 507374 -284
rect 507430 -340 507498 -284
rect 507554 -340 507622 -284
rect 507678 -340 507774 -284
rect 507154 -408 507774 -340
rect 507154 -464 507250 -408
rect 507306 -464 507374 -408
rect 507430 -464 507498 -408
rect 507554 -464 507622 -408
rect 507678 -464 507774 -408
rect 507154 -532 507774 -464
rect 507154 -588 507250 -532
rect 507306 -588 507374 -532
rect 507430 -588 507498 -532
rect 507554 -588 507622 -532
rect 507678 -588 507774 -532
rect 507154 -1644 507774 -588
rect 510874 28350 511494 32890
rect 510874 28294 510970 28350
rect 511026 28294 511094 28350
rect 511150 28294 511218 28350
rect 511274 28294 511342 28350
rect 511398 28294 511494 28350
rect 510874 28226 511494 28294
rect 510874 28170 510970 28226
rect 511026 28170 511094 28226
rect 511150 28170 511218 28226
rect 511274 28170 511342 28226
rect 511398 28170 511494 28226
rect 510874 28102 511494 28170
rect 510874 28046 510970 28102
rect 511026 28046 511094 28102
rect 511150 28046 511218 28102
rect 511274 28046 511342 28102
rect 511398 28046 511494 28102
rect 510874 27978 511494 28046
rect 510874 27922 510970 27978
rect 511026 27922 511094 27978
rect 511150 27922 511218 27978
rect 511274 27922 511342 27978
rect 511398 27922 511494 27978
rect 510874 10350 511494 27922
rect 510874 10294 510970 10350
rect 511026 10294 511094 10350
rect 511150 10294 511218 10350
rect 511274 10294 511342 10350
rect 511398 10294 511494 10350
rect 510874 10226 511494 10294
rect 510874 10170 510970 10226
rect 511026 10170 511094 10226
rect 511150 10170 511218 10226
rect 511274 10170 511342 10226
rect 511398 10170 511494 10226
rect 510874 10102 511494 10170
rect 510874 10046 510970 10102
rect 511026 10046 511094 10102
rect 511150 10046 511218 10102
rect 511274 10046 511342 10102
rect 511398 10046 511494 10102
rect 510874 9978 511494 10046
rect 510874 9922 510970 9978
rect 511026 9922 511094 9978
rect 511150 9922 511218 9978
rect 511274 9922 511342 9978
rect 511398 9922 511494 9978
rect 510874 -1120 511494 9922
rect 510874 -1176 510970 -1120
rect 511026 -1176 511094 -1120
rect 511150 -1176 511218 -1120
rect 511274 -1176 511342 -1120
rect 511398 -1176 511494 -1120
rect 510874 -1244 511494 -1176
rect 510874 -1300 510970 -1244
rect 511026 -1300 511094 -1244
rect 511150 -1300 511218 -1244
rect 511274 -1300 511342 -1244
rect 511398 -1300 511494 -1244
rect 510874 -1368 511494 -1300
rect 510874 -1424 510970 -1368
rect 511026 -1424 511094 -1368
rect 511150 -1424 511218 -1368
rect 511274 -1424 511342 -1368
rect 511398 -1424 511494 -1368
rect 510874 -1492 511494 -1424
rect 510874 -1548 510970 -1492
rect 511026 -1548 511094 -1492
rect 511150 -1548 511218 -1492
rect 511274 -1548 511342 -1492
rect 511398 -1548 511494 -1492
rect 510874 -1644 511494 -1548
rect 525154 22350 525774 32890
rect 525154 22294 525250 22350
rect 525306 22294 525374 22350
rect 525430 22294 525498 22350
rect 525554 22294 525622 22350
rect 525678 22294 525774 22350
rect 525154 22226 525774 22294
rect 525154 22170 525250 22226
rect 525306 22170 525374 22226
rect 525430 22170 525498 22226
rect 525554 22170 525622 22226
rect 525678 22170 525774 22226
rect 525154 22102 525774 22170
rect 525154 22046 525250 22102
rect 525306 22046 525374 22102
rect 525430 22046 525498 22102
rect 525554 22046 525622 22102
rect 525678 22046 525774 22102
rect 525154 21978 525774 22046
rect 525154 21922 525250 21978
rect 525306 21922 525374 21978
rect 525430 21922 525498 21978
rect 525554 21922 525622 21978
rect 525678 21922 525774 21978
rect 525154 4350 525774 21922
rect 525154 4294 525250 4350
rect 525306 4294 525374 4350
rect 525430 4294 525498 4350
rect 525554 4294 525622 4350
rect 525678 4294 525774 4350
rect 525154 4226 525774 4294
rect 525154 4170 525250 4226
rect 525306 4170 525374 4226
rect 525430 4170 525498 4226
rect 525554 4170 525622 4226
rect 525678 4170 525774 4226
rect 525154 4102 525774 4170
rect 525154 4046 525250 4102
rect 525306 4046 525374 4102
rect 525430 4046 525498 4102
rect 525554 4046 525622 4102
rect 525678 4046 525774 4102
rect 525154 3978 525774 4046
rect 525154 3922 525250 3978
rect 525306 3922 525374 3978
rect 525430 3922 525498 3978
rect 525554 3922 525622 3978
rect 525678 3922 525774 3978
rect 525154 -160 525774 3922
rect 525154 -216 525250 -160
rect 525306 -216 525374 -160
rect 525430 -216 525498 -160
rect 525554 -216 525622 -160
rect 525678 -216 525774 -160
rect 525154 -284 525774 -216
rect 525154 -340 525250 -284
rect 525306 -340 525374 -284
rect 525430 -340 525498 -284
rect 525554 -340 525622 -284
rect 525678 -340 525774 -284
rect 525154 -408 525774 -340
rect 525154 -464 525250 -408
rect 525306 -464 525374 -408
rect 525430 -464 525498 -408
rect 525554 -464 525622 -408
rect 525678 -464 525774 -408
rect 525154 -532 525774 -464
rect 525154 -588 525250 -532
rect 525306 -588 525374 -532
rect 525430 -588 525498 -532
rect 525554 -588 525622 -532
rect 525678 -588 525774 -532
rect 525154 -1644 525774 -588
rect 528874 28350 529494 32890
rect 528874 28294 528970 28350
rect 529026 28294 529094 28350
rect 529150 28294 529218 28350
rect 529274 28294 529342 28350
rect 529398 28294 529494 28350
rect 528874 28226 529494 28294
rect 528874 28170 528970 28226
rect 529026 28170 529094 28226
rect 529150 28170 529218 28226
rect 529274 28170 529342 28226
rect 529398 28170 529494 28226
rect 528874 28102 529494 28170
rect 528874 28046 528970 28102
rect 529026 28046 529094 28102
rect 529150 28046 529218 28102
rect 529274 28046 529342 28102
rect 529398 28046 529494 28102
rect 528874 27978 529494 28046
rect 528874 27922 528970 27978
rect 529026 27922 529094 27978
rect 529150 27922 529218 27978
rect 529274 27922 529342 27978
rect 529398 27922 529494 27978
rect 528874 10350 529494 27922
rect 528874 10294 528970 10350
rect 529026 10294 529094 10350
rect 529150 10294 529218 10350
rect 529274 10294 529342 10350
rect 529398 10294 529494 10350
rect 528874 10226 529494 10294
rect 528874 10170 528970 10226
rect 529026 10170 529094 10226
rect 529150 10170 529218 10226
rect 529274 10170 529342 10226
rect 529398 10170 529494 10226
rect 528874 10102 529494 10170
rect 528874 10046 528970 10102
rect 529026 10046 529094 10102
rect 529150 10046 529218 10102
rect 529274 10046 529342 10102
rect 529398 10046 529494 10102
rect 528874 9978 529494 10046
rect 528874 9922 528970 9978
rect 529026 9922 529094 9978
rect 529150 9922 529218 9978
rect 529274 9922 529342 9978
rect 529398 9922 529494 9978
rect 528874 -1120 529494 9922
rect 528874 -1176 528970 -1120
rect 529026 -1176 529094 -1120
rect 529150 -1176 529218 -1120
rect 529274 -1176 529342 -1120
rect 529398 -1176 529494 -1120
rect 528874 -1244 529494 -1176
rect 528874 -1300 528970 -1244
rect 529026 -1300 529094 -1244
rect 529150 -1300 529218 -1244
rect 529274 -1300 529342 -1244
rect 529398 -1300 529494 -1244
rect 528874 -1368 529494 -1300
rect 528874 -1424 528970 -1368
rect 529026 -1424 529094 -1368
rect 529150 -1424 529218 -1368
rect 529274 -1424 529342 -1368
rect 529398 -1424 529494 -1368
rect 528874 -1492 529494 -1424
rect 528874 -1548 528970 -1492
rect 529026 -1548 529094 -1492
rect 529150 -1548 529218 -1492
rect 529274 -1548 529342 -1492
rect 529398 -1548 529494 -1492
rect 528874 -1644 529494 -1548
rect 543154 22350 543774 32890
rect 543154 22294 543250 22350
rect 543306 22294 543374 22350
rect 543430 22294 543498 22350
rect 543554 22294 543622 22350
rect 543678 22294 543774 22350
rect 543154 22226 543774 22294
rect 543154 22170 543250 22226
rect 543306 22170 543374 22226
rect 543430 22170 543498 22226
rect 543554 22170 543622 22226
rect 543678 22170 543774 22226
rect 543154 22102 543774 22170
rect 543154 22046 543250 22102
rect 543306 22046 543374 22102
rect 543430 22046 543498 22102
rect 543554 22046 543622 22102
rect 543678 22046 543774 22102
rect 543154 21978 543774 22046
rect 543154 21922 543250 21978
rect 543306 21922 543374 21978
rect 543430 21922 543498 21978
rect 543554 21922 543622 21978
rect 543678 21922 543774 21978
rect 543154 4350 543774 21922
rect 543154 4294 543250 4350
rect 543306 4294 543374 4350
rect 543430 4294 543498 4350
rect 543554 4294 543622 4350
rect 543678 4294 543774 4350
rect 543154 4226 543774 4294
rect 543154 4170 543250 4226
rect 543306 4170 543374 4226
rect 543430 4170 543498 4226
rect 543554 4170 543622 4226
rect 543678 4170 543774 4226
rect 543154 4102 543774 4170
rect 543154 4046 543250 4102
rect 543306 4046 543374 4102
rect 543430 4046 543498 4102
rect 543554 4046 543622 4102
rect 543678 4046 543774 4102
rect 543154 3978 543774 4046
rect 543154 3922 543250 3978
rect 543306 3922 543374 3978
rect 543430 3922 543498 3978
rect 543554 3922 543622 3978
rect 543678 3922 543774 3978
rect 543154 -160 543774 3922
rect 543154 -216 543250 -160
rect 543306 -216 543374 -160
rect 543430 -216 543498 -160
rect 543554 -216 543622 -160
rect 543678 -216 543774 -160
rect 543154 -284 543774 -216
rect 543154 -340 543250 -284
rect 543306 -340 543374 -284
rect 543430 -340 543498 -284
rect 543554 -340 543622 -284
rect 543678 -340 543774 -284
rect 543154 -408 543774 -340
rect 543154 -464 543250 -408
rect 543306 -464 543374 -408
rect 543430 -464 543498 -408
rect 543554 -464 543622 -408
rect 543678 -464 543774 -408
rect 543154 -532 543774 -464
rect 543154 -588 543250 -532
rect 543306 -588 543374 -532
rect 543430 -588 543498 -532
rect 543554 -588 543622 -532
rect 543678 -588 543774 -532
rect 543154 -1644 543774 -588
rect 546874 28350 547494 32890
rect 546874 28294 546970 28350
rect 547026 28294 547094 28350
rect 547150 28294 547218 28350
rect 547274 28294 547342 28350
rect 547398 28294 547494 28350
rect 546874 28226 547494 28294
rect 546874 28170 546970 28226
rect 547026 28170 547094 28226
rect 547150 28170 547218 28226
rect 547274 28170 547342 28226
rect 547398 28170 547494 28226
rect 546874 28102 547494 28170
rect 546874 28046 546970 28102
rect 547026 28046 547094 28102
rect 547150 28046 547218 28102
rect 547274 28046 547342 28102
rect 547398 28046 547494 28102
rect 546874 27978 547494 28046
rect 546874 27922 546970 27978
rect 547026 27922 547094 27978
rect 547150 27922 547218 27978
rect 547274 27922 547342 27978
rect 547398 27922 547494 27978
rect 546874 10350 547494 27922
rect 546874 10294 546970 10350
rect 547026 10294 547094 10350
rect 547150 10294 547218 10350
rect 547274 10294 547342 10350
rect 547398 10294 547494 10350
rect 546874 10226 547494 10294
rect 546874 10170 546970 10226
rect 547026 10170 547094 10226
rect 547150 10170 547218 10226
rect 547274 10170 547342 10226
rect 547398 10170 547494 10226
rect 546874 10102 547494 10170
rect 546874 10046 546970 10102
rect 547026 10046 547094 10102
rect 547150 10046 547218 10102
rect 547274 10046 547342 10102
rect 547398 10046 547494 10102
rect 546874 9978 547494 10046
rect 546874 9922 546970 9978
rect 547026 9922 547094 9978
rect 547150 9922 547218 9978
rect 547274 9922 547342 9978
rect 547398 9922 547494 9978
rect 546874 -1120 547494 9922
rect 546874 -1176 546970 -1120
rect 547026 -1176 547094 -1120
rect 547150 -1176 547218 -1120
rect 547274 -1176 547342 -1120
rect 547398 -1176 547494 -1120
rect 546874 -1244 547494 -1176
rect 546874 -1300 546970 -1244
rect 547026 -1300 547094 -1244
rect 547150 -1300 547218 -1244
rect 547274 -1300 547342 -1244
rect 547398 -1300 547494 -1244
rect 546874 -1368 547494 -1300
rect 546874 -1424 546970 -1368
rect 547026 -1424 547094 -1368
rect 547150 -1424 547218 -1368
rect 547274 -1424 547342 -1368
rect 547398 -1424 547494 -1368
rect 546874 -1492 547494 -1424
rect 546874 -1548 546970 -1492
rect 547026 -1548 547094 -1492
rect 547150 -1548 547218 -1492
rect 547274 -1548 547342 -1492
rect 547398 -1548 547494 -1492
rect 546874 -1644 547494 -1548
rect 561154 22350 561774 39922
rect 561154 22294 561250 22350
rect 561306 22294 561374 22350
rect 561430 22294 561498 22350
rect 561554 22294 561622 22350
rect 561678 22294 561774 22350
rect 561154 22226 561774 22294
rect 561154 22170 561250 22226
rect 561306 22170 561374 22226
rect 561430 22170 561498 22226
rect 561554 22170 561622 22226
rect 561678 22170 561774 22226
rect 561154 22102 561774 22170
rect 561154 22046 561250 22102
rect 561306 22046 561374 22102
rect 561430 22046 561498 22102
rect 561554 22046 561622 22102
rect 561678 22046 561774 22102
rect 561154 21978 561774 22046
rect 561154 21922 561250 21978
rect 561306 21922 561374 21978
rect 561430 21922 561498 21978
rect 561554 21922 561622 21978
rect 561678 21922 561774 21978
rect 561154 4350 561774 21922
rect 561154 4294 561250 4350
rect 561306 4294 561374 4350
rect 561430 4294 561498 4350
rect 561554 4294 561622 4350
rect 561678 4294 561774 4350
rect 561154 4226 561774 4294
rect 561154 4170 561250 4226
rect 561306 4170 561374 4226
rect 561430 4170 561498 4226
rect 561554 4170 561622 4226
rect 561678 4170 561774 4226
rect 561154 4102 561774 4170
rect 561154 4046 561250 4102
rect 561306 4046 561374 4102
rect 561430 4046 561498 4102
rect 561554 4046 561622 4102
rect 561678 4046 561774 4102
rect 561154 3978 561774 4046
rect 561154 3922 561250 3978
rect 561306 3922 561374 3978
rect 561430 3922 561498 3978
rect 561554 3922 561622 3978
rect 561678 3922 561774 3978
rect 561154 -160 561774 3922
rect 561154 -216 561250 -160
rect 561306 -216 561374 -160
rect 561430 -216 561498 -160
rect 561554 -216 561622 -160
rect 561678 -216 561774 -160
rect 561154 -284 561774 -216
rect 561154 -340 561250 -284
rect 561306 -340 561374 -284
rect 561430 -340 561498 -284
rect 561554 -340 561622 -284
rect 561678 -340 561774 -284
rect 561154 -408 561774 -340
rect 561154 -464 561250 -408
rect 561306 -464 561374 -408
rect 561430 -464 561498 -408
rect 561554 -464 561622 -408
rect 561678 -464 561774 -408
rect 561154 -532 561774 -464
rect 561154 -588 561250 -532
rect 561306 -588 561374 -532
rect 561430 -588 561498 -532
rect 561554 -588 561622 -532
rect 561678 -588 561774 -532
rect 561154 -1644 561774 -588
rect 564874 598172 565494 598268
rect 564874 598116 564970 598172
rect 565026 598116 565094 598172
rect 565150 598116 565218 598172
rect 565274 598116 565342 598172
rect 565398 598116 565494 598172
rect 564874 598048 565494 598116
rect 564874 597992 564970 598048
rect 565026 597992 565094 598048
rect 565150 597992 565218 598048
rect 565274 597992 565342 598048
rect 565398 597992 565494 598048
rect 564874 597924 565494 597992
rect 564874 597868 564970 597924
rect 565026 597868 565094 597924
rect 565150 597868 565218 597924
rect 565274 597868 565342 597924
rect 565398 597868 565494 597924
rect 564874 597800 565494 597868
rect 564874 597744 564970 597800
rect 565026 597744 565094 597800
rect 565150 597744 565218 597800
rect 565274 597744 565342 597800
rect 565398 597744 565494 597800
rect 564874 586350 565494 597744
rect 564874 586294 564970 586350
rect 565026 586294 565094 586350
rect 565150 586294 565218 586350
rect 565274 586294 565342 586350
rect 565398 586294 565494 586350
rect 564874 586226 565494 586294
rect 564874 586170 564970 586226
rect 565026 586170 565094 586226
rect 565150 586170 565218 586226
rect 565274 586170 565342 586226
rect 565398 586170 565494 586226
rect 564874 586102 565494 586170
rect 564874 586046 564970 586102
rect 565026 586046 565094 586102
rect 565150 586046 565218 586102
rect 565274 586046 565342 586102
rect 565398 586046 565494 586102
rect 564874 585978 565494 586046
rect 564874 585922 564970 585978
rect 565026 585922 565094 585978
rect 565150 585922 565218 585978
rect 565274 585922 565342 585978
rect 565398 585922 565494 585978
rect 564874 568350 565494 585922
rect 564874 568294 564970 568350
rect 565026 568294 565094 568350
rect 565150 568294 565218 568350
rect 565274 568294 565342 568350
rect 565398 568294 565494 568350
rect 564874 568226 565494 568294
rect 564874 568170 564970 568226
rect 565026 568170 565094 568226
rect 565150 568170 565218 568226
rect 565274 568170 565342 568226
rect 565398 568170 565494 568226
rect 564874 568102 565494 568170
rect 564874 568046 564970 568102
rect 565026 568046 565094 568102
rect 565150 568046 565218 568102
rect 565274 568046 565342 568102
rect 565398 568046 565494 568102
rect 564874 567978 565494 568046
rect 564874 567922 564970 567978
rect 565026 567922 565094 567978
rect 565150 567922 565218 567978
rect 565274 567922 565342 567978
rect 565398 567922 565494 567978
rect 564874 550350 565494 567922
rect 564874 550294 564970 550350
rect 565026 550294 565094 550350
rect 565150 550294 565218 550350
rect 565274 550294 565342 550350
rect 565398 550294 565494 550350
rect 564874 550226 565494 550294
rect 564874 550170 564970 550226
rect 565026 550170 565094 550226
rect 565150 550170 565218 550226
rect 565274 550170 565342 550226
rect 565398 550170 565494 550226
rect 564874 550102 565494 550170
rect 564874 550046 564970 550102
rect 565026 550046 565094 550102
rect 565150 550046 565218 550102
rect 565274 550046 565342 550102
rect 565398 550046 565494 550102
rect 564874 549978 565494 550046
rect 564874 549922 564970 549978
rect 565026 549922 565094 549978
rect 565150 549922 565218 549978
rect 565274 549922 565342 549978
rect 565398 549922 565494 549978
rect 564874 532350 565494 549922
rect 564874 532294 564970 532350
rect 565026 532294 565094 532350
rect 565150 532294 565218 532350
rect 565274 532294 565342 532350
rect 565398 532294 565494 532350
rect 564874 532226 565494 532294
rect 564874 532170 564970 532226
rect 565026 532170 565094 532226
rect 565150 532170 565218 532226
rect 565274 532170 565342 532226
rect 565398 532170 565494 532226
rect 564874 532102 565494 532170
rect 564874 532046 564970 532102
rect 565026 532046 565094 532102
rect 565150 532046 565218 532102
rect 565274 532046 565342 532102
rect 565398 532046 565494 532102
rect 564874 531978 565494 532046
rect 564874 531922 564970 531978
rect 565026 531922 565094 531978
rect 565150 531922 565218 531978
rect 565274 531922 565342 531978
rect 565398 531922 565494 531978
rect 564874 514350 565494 531922
rect 564874 514294 564970 514350
rect 565026 514294 565094 514350
rect 565150 514294 565218 514350
rect 565274 514294 565342 514350
rect 565398 514294 565494 514350
rect 564874 514226 565494 514294
rect 564874 514170 564970 514226
rect 565026 514170 565094 514226
rect 565150 514170 565218 514226
rect 565274 514170 565342 514226
rect 565398 514170 565494 514226
rect 564874 514102 565494 514170
rect 564874 514046 564970 514102
rect 565026 514046 565094 514102
rect 565150 514046 565218 514102
rect 565274 514046 565342 514102
rect 565398 514046 565494 514102
rect 564874 513978 565494 514046
rect 564874 513922 564970 513978
rect 565026 513922 565094 513978
rect 565150 513922 565218 513978
rect 565274 513922 565342 513978
rect 565398 513922 565494 513978
rect 564874 496350 565494 513922
rect 564874 496294 564970 496350
rect 565026 496294 565094 496350
rect 565150 496294 565218 496350
rect 565274 496294 565342 496350
rect 565398 496294 565494 496350
rect 564874 496226 565494 496294
rect 564874 496170 564970 496226
rect 565026 496170 565094 496226
rect 565150 496170 565218 496226
rect 565274 496170 565342 496226
rect 565398 496170 565494 496226
rect 564874 496102 565494 496170
rect 564874 496046 564970 496102
rect 565026 496046 565094 496102
rect 565150 496046 565218 496102
rect 565274 496046 565342 496102
rect 565398 496046 565494 496102
rect 564874 495978 565494 496046
rect 564874 495922 564970 495978
rect 565026 495922 565094 495978
rect 565150 495922 565218 495978
rect 565274 495922 565342 495978
rect 565398 495922 565494 495978
rect 564874 478350 565494 495922
rect 564874 478294 564970 478350
rect 565026 478294 565094 478350
rect 565150 478294 565218 478350
rect 565274 478294 565342 478350
rect 565398 478294 565494 478350
rect 564874 478226 565494 478294
rect 564874 478170 564970 478226
rect 565026 478170 565094 478226
rect 565150 478170 565218 478226
rect 565274 478170 565342 478226
rect 565398 478170 565494 478226
rect 564874 478102 565494 478170
rect 564874 478046 564970 478102
rect 565026 478046 565094 478102
rect 565150 478046 565218 478102
rect 565274 478046 565342 478102
rect 565398 478046 565494 478102
rect 564874 477978 565494 478046
rect 564874 477922 564970 477978
rect 565026 477922 565094 477978
rect 565150 477922 565218 477978
rect 565274 477922 565342 477978
rect 565398 477922 565494 477978
rect 564874 460350 565494 477922
rect 564874 460294 564970 460350
rect 565026 460294 565094 460350
rect 565150 460294 565218 460350
rect 565274 460294 565342 460350
rect 565398 460294 565494 460350
rect 564874 460226 565494 460294
rect 564874 460170 564970 460226
rect 565026 460170 565094 460226
rect 565150 460170 565218 460226
rect 565274 460170 565342 460226
rect 565398 460170 565494 460226
rect 564874 460102 565494 460170
rect 564874 460046 564970 460102
rect 565026 460046 565094 460102
rect 565150 460046 565218 460102
rect 565274 460046 565342 460102
rect 565398 460046 565494 460102
rect 564874 459978 565494 460046
rect 564874 459922 564970 459978
rect 565026 459922 565094 459978
rect 565150 459922 565218 459978
rect 565274 459922 565342 459978
rect 565398 459922 565494 459978
rect 564874 442350 565494 459922
rect 564874 442294 564970 442350
rect 565026 442294 565094 442350
rect 565150 442294 565218 442350
rect 565274 442294 565342 442350
rect 565398 442294 565494 442350
rect 564874 442226 565494 442294
rect 564874 442170 564970 442226
rect 565026 442170 565094 442226
rect 565150 442170 565218 442226
rect 565274 442170 565342 442226
rect 565398 442170 565494 442226
rect 564874 442102 565494 442170
rect 564874 442046 564970 442102
rect 565026 442046 565094 442102
rect 565150 442046 565218 442102
rect 565274 442046 565342 442102
rect 565398 442046 565494 442102
rect 564874 441978 565494 442046
rect 564874 441922 564970 441978
rect 565026 441922 565094 441978
rect 565150 441922 565218 441978
rect 565274 441922 565342 441978
rect 565398 441922 565494 441978
rect 564874 424350 565494 441922
rect 564874 424294 564970 424350
rect 565026 424294 565094 424350
rect 565150 424294 565218 424350
rect 565274 424294 565342 424350
rect 565398 424294 565494 424350
rect 564874 424226 565494 424294
rect 564874 424170 564970 424226
rect 565026 424170 565094 424226
rect 565150 424170 565218 424226
rect 565274 424170 565342 424226
rect 565398 424170 565494 424226
rect 564874 424102 565494 424170
rect 564874 424046 564970 424102
rect 565026 424046 565094 424102
rect 565150 424046 565218 424102
rect 565274 424046 565342 424102
rect 565398 424046 565494 424102
rect 564874 423978 565494 424046
rect 564874 423922 564970 423978
rect 565026 423922 565094 423978
rect 565150 423922 565218 423978
rect 565274 423922 565342 423978
rect 565398 423922 565494 423978
rect 564874 406350 565494 423922
rect 564874 406294 564970 406350
rect 565026 406294 565094 406350
rect 565150 406294 565218 406350
rect 565274 406294 565342 406350
rect 565398 406294 565494 406350
rect 564874 406226 565494 406294
rect 564874 406170 564970 406226
rect 565026 406170 565094 406226
rect 565150 406170 565218 406226
rect 565274 406170 565342 406226
rect 565398 406170 565494 406226
rect 564874 406102 565494 406170
rect 564874 406046 564970 406102
rect 565026 406046 565094 406102
rect 565150 406046 565218 406102
rect 565274 406046 565342 406102
rect 565398 406046 565494 406102
rect 564874 405978 565494 406046
rect 564874 405922 564970 405978
rect 565026 405922 565094 405978
rect 565150 405922 565218 405978
rect 565274 405922 565342 405978
rect 565398 405922 565494 405978
rect 564874 388350 565494 405922
rect 564874 388294 564970 388350
rect 565026 388294 565094 388350
rect 565150 388294 565218 388350
rect 565274 388294 565342 388350
rect 565398 388294 565494 388350
rect 564874 388226 565494 388294
rect 564874 388170 564970 388226
rect 565026 388170 565094 388226
rect 565150 388170 565218 388226
rect 565274 388170 565342 388226
rect 565398 388170 565494 388226
rect 564874 388102 565494 388170
rect 564874 388046 564970 388102
rect 565026 388046 565094 388102
rect 565150 388046 565218 388102
rect 565274 388046 565342 388102
rect 565398 388046 565494 388102
rect 564874 387978 565494 388046
rect 564874 387922 564970 387978
rect 565026 387922 565094 387978
rect 565150 387922 565218 387978
rect 565274 387922 565342 387978
rect 565398 387922 565494 387978
rect 564874 370350 565494 387922
rect 564874 370294 564970 370350
rect 565026 370294 565094 370350
rect 565150 370294 565218 370350
rect 565274 370294 565342 370350
rect 565398 370294 565494 370350
rect 564874 370226 565494 370294
rect 564874 370170 564970 370226
rect 565026 370170 565094 370226
rect 565150 370170 565218 370226
rect 565274 370170 565342 370226
rect 565398 370170 565494 370226
rect 564874 370102 565494 370170
rect 564874 370046 564970 370102
rect 565026 370046 565094 370102
rect 565150 370046 565218 370102
rect 565274 370046 565342 370102
rect 565398 370046 565494 370102
rect 564874 369978 565494 370046
rect 564874 369922 564970 369978
rect 565026 369922 565094 369978
rect 565150 369922 565218 369978
rect 565274 369922 565342 369978
rect 565398 369922 565494 369978
rect 564874 352350 565494 369922
rect 564874 352294 564970 352350
rect 565026 352294 565094 352350
rect 565150 352294 565218 352350
rect 565274 352294 565342 352350
rect 565398 352294 565494 352350
rect 564874 352226 565494 352294
rect 564874 352170 564970 352226
rect 565026 352170 565094 352226
rect 565150 352170 565218 352226
rect 565274 352170 565342 352226
rect 565398 352170 565494 352226
rect 564874 352102 565494 352170
rect 564874 352046 564970 352102
rect 565026 352046 565094 352102
rect 565150 352046 565218 352102
rect 565274 352046 565342 352102
rect 565398 352046 565494 352102
rect 564874 351978 565494 352046
rect 564874 351922 564970 351978
rect 565026 351922 565094 351978
rect 565150 351922 565218 351978
rect 565274 351922 565342 351978
rect 565398 351922 565494 351978
rect 564874 334350 565494 351922
rect 564874 334294 564970 334350
rect 565026 334294 565094 334350
rect 565150 334294 565218 334350
rect 565274 334294 565342 334350
rect 565398 334294 565494 334350
rect 564874 334226 565494 334294
rect 564874 334170 564970 334226
rect 565026 334170 565094 334226
rect 565150 334170 565218 334226
rect 565274 334170 565342 334226
rect 565398 334170 565494 334226
rect 564874 334102 565494 334170
rect 564874 334046 564970 334102
rect 565026 334046 565094 334102
rect 565150 334046 565218 334102
rect 565274 334046 565342 334102
rect 565398 334046 565494 334102
rect 564874 333978 565494 334046
rect 564874 333922 564970 333978
rect 565026 333922 565094 333978
rect 565150 333922 565218 333978
rect 565274 333922 565342 333978
rect 565398 333922 565494 333978
rect 564874 316350 565494 333922
rect 564874 316294 564970 316350
rect 565026 316294 565094 316350
rect 565150 316294 565218 316350
rect 565274 316294 565342 316350
rect 565398 316294 565494 316350
rect 564874 316226 565494 316294
rect 564874 316170 564970 316226
rect 565026 316170 565094 316226
rect 565150 316170 565218 316226
rect 565274 316170 565342 316226
rect 565398 316170 565494 316226
rect 564874 316102 565494 316170
rect 564874 316046 564970 316102
rect 565026 316046 565094 316102
rect 565150 316046 565218 316102
rect 565274 316046 565342 316102
rect 565398 316046 565494 316102
rect 564874 315978 565494 316046
rect 564874 315922 564970 315978
rect 565026 315922 565094 315978
rect 565150 315922 565218 315978
rect 565274 315922 565342 315978
rect 565398 315922 565494 315978
rect 564874 298350 565494 315922
rect 564874 298294 564970 298350
rect 565026 298294 565094 298350
rect 565150 298294 565218 298350
rect 565274 298294 565342 298350
rect 565398 298294 565494 298350
rect 564874 298226 565494 298294
rect 564874 298170 564970 298226
rect 565026 298170 565094 298226
rect 565150 298170 565218 298226
rect 565274 298170 565342 298226
rect 565398 298170 565494 298226
rect 564874 298102 565494 298170
rect 564874 298046 564970 298102
rect 565026 298046 565094 298102
rect 565150 298046 565218 298102
rect 565274 298046 565342 298102
rect 565398 298046 565494 298102
rect 564874 297978 565494 298046
rect 564874 297922 564970 297978
rect 565026 297922 565094 297978
rect 565150 297922 565218 297978
rect 565274 297922 565342 297978
rect 565398 297922 565494 297978
rect 564874 280350 565494 297922
rect 564874 280294 564970 280350
rect 565026 280294 565094 280350
rect 565150 280294 565218 280350
rect 565274 280294 565342 280350
rect 565398 280294 565494 280350
rect 564874 280226 565494 280294
rect 564874 280170 564970 280226
rect 565026 280170 565094 280226
rect 565150 280170 565218 280226
rect 565274 280170 565342 280226
rect 565398 280170 565494 280226
rect 564874 280102 565494 280170
rect 564874 280046 564970 280102
rect 565026 280046 565094 280102
rect 565150 280046 565218 280102
rect 565274 280046 565342 280102
rect 565398 280046 565494 280102
rect 564874 279978 565494 280046
rect 564874 279922 564970 279978
rect 565026 279922 565094 279978
rect 565150 279922 565218 279978
rect 565274 279922 565342 279978
rect 565398 279922 565494 279978
rect 564874 262350 565494 279922
rect 564874 262294 564970 262350
rect 565026 262294 565094 262350
rect 565150 262294 565218 262350
rect 565274 262294 565342 262350
rect 565398 262294 565494 262350
rect 564874 262226 565494 262294
rect 564874 262170 564970 262226
rect 565026 262170 565094 262226
rect 565150 262170 565218 262226
rect 565274 262170 565342 262226
rect 565398 262170 565494 262226
rect 564874 262102 565494 262170
rect 564874 262046 564970 262102
rect 565026 262046 565094 262102
rect 565150 262046 565218 262102
rect 565274 262046 565342 262102
rect 565398 262046 565494 262102
rect 564874 261978 565494 262046
rect 564874 261922 564970 261978
rect 565026 261922 565094 261978
rect 565150 261922 565218 261978
rect 565274 261922 565342 261978
rect 565398 261922 565494 261978
rect 564874 244350 565494 261922
rect 564874 244294 564970 244350
rect 565026 244294 565094 244350
rect 565150 244294 565218 244350
rect 565274 244294 565342 244350
rect 565398 244294 565494 244350
rect 564874 244226 565494 244294
rect 564874 244170 564970 244226
rect 565026 244170 565094 244226
rect 565150 244170 565218 244226
rect 565274 244170 565342 244226
rect 565398 244170 565494 244226
rect 564874 244102 565494 244170
rect 564874 244046 564970 244102
rect 565026 244046 565094 244102
rect 565150 244046 565218 244102
rect 565274 244046 565342 244102
rect 565398 244046 565494 244102
rect 564874 243978 565494 244046
rect 564874 243922 564970 243978
rect 565026 243922 565094 243978
rect 565150 243922 565218 243978
rect 565274 243922 565342 243978
rect 565398 243922 565494 243978
rect 564874 226350 565494 243922
rect 564874 226294 564970 226350
rect 565026 226294 565094 226350
rect 565150 226294 565218 226350
rect 565274 226294 565342 226350
rect 565398 226294 565494 226350
rect 564874 226226 565494 226294
rect 564874 226170 564970 226226
rect 565026 226170 565094 226226
rect 565150 226170 565218 226226
rect 565274 226170 565342 226226
rect 565398 226170 565494 226226
rect 564874 226102 565494 226170
rect 564874 226046 564970 226102
rect 565026 226046 565094 226102
rect 565150 226046 565218 226102
rect 565274 226046 565342 226102
rect 565398 226046 565494 226102
rect 564874 225978 565494 226046
rect 564874 225922 564970 225978
rect 565026 225922 565094 225978
rect 565150 225922 565218 225978
rect 565274 225922 565342 225978
rect 565398 225922 565494 225978
rect 564874 208350 565494 225922
rect 564874 208294 564970 208350
rect 565026 208294 565094 208350
rect 565150 208294 565218 208350
rect 565274 208294 565342 208350
rect 565398 208294 565494 208350
rect 564874 208226 565494 208294
rect 564874 208170 564970 208226
rect 565026 208170 565094 208226
rect 565150 208170 565218 208226
rect 565274 208170 565342 208226
rect 565398 208170 565494 208226
rect 564874 208102 565494 208170
rect 564874 208046 564970 208102
rect 565026 208046 565094 208102
rect 565150 208046 565218 208102
rect 565274 208046 565342 208102
rect 565398 208046 565494 208102
rect 564874 207978 565494 208046
rect 564874 207922 564970 207978
rect 565026 207922 565094 207978
rect 565150 207922 565218 207978
rect 565274 207922 565342 207978
rect 565398 207922 565494 207978
rect 564874 190350 565494 207922
rect 564874 190294 564970 190350
rect 565026 190294 565094 190350
rect 565150 190294 565218 190350
rect 565274 190294 565342 190350
rect 565398 190294 565494 190350
rect 564874 190226 565494 190294
rect 564874 190170 564970 190226
rect 565026 190170 565094 190226
rect 565150 190170 565218 190226
rect 565274 190170 565342 190226
rect 565398 190170 565494 190226
rect 564874 190102 565494 190170
rect 564874 190046 564970 190102
rect 565026 190046 565094 190102
rect 565150 190046 565218 190102
rect 565274 190046 565342 190102
rect 565398 190046 565494 190102
rect 564874 189978 565494 190046
rect 564874 189922 564970 189978
rect 565026 189922 565094 189978
rect 565150 189922 565218 189978
rect 565274 189922 565342 189978
rect 565398 189922 565494 189978
rect 564874 172350 565494 189922
rect 564874 172294 564970 172350
rect 565026 172294 565094 172350
rect 565150 172294 565218 172350
rect 565274 172294 565342 172350
rect 565398 172294 565494 172350
rect 564874 172226 565494 172294
rect 564874 172170 564970 172226
rect 565026 172170 565094 172226
rect 565150 172170 565218 172226
rect 565274 172170 565342 172226
rect 565398 172170 565494 172226
rect 564874 172102 565494 172170
rect 564874 172046 564970 172102
rect 565026 172046 565094 172102
rect 565150 172046 565218 172102
rect 565274 172046 565342 172102
rect 565398 172046 565494 172102
rect 564874 171978 565494 172046
rect 564874 171922 564970 171978
rect 565026 171922 565094 171978
rect 565150 171922 565218 171978
rect 565274 171922 565342 171978
rect 565398 171922 565494 171978
rect 564874 154350 565494 171922
rect 564874 154294 564970 154350
rect 565026 154294 565094 154350
rect 565150 154294 565218 154350
rect 565274 154294 565342 154350
rect 565398 154294 565494 154350
rect 564874 154226 565494 154294
rect 564874 154170 564970 154226
rect 565026 154170 565094 154226
rect 565150 154170 565218 154226
rect 565274 154170 565342 154226
rect 565398 154170 565494 154226
rect 564874 154102 565494 154170
rect 564874 154046 564970 154102
rect 565026 154046 565094 154102
rect 565150 154046 565218 154102
rect 565274 154046 565342 154102
rect 565398 154046 565494 154102
rect 564874 153978 565494 154046
rect 564874 153922 564970 153978
rect 565026 153922 565094 153978
rect 565150 153922 565218 153978
rect 565274 153922 565342 153978
rect 565398 153922 565494 153978
rect 564874 136350 565494 153922
rect 564874 136294 564970 136350
rect 565026 136294 565094 136350
rect 565150 136294 565218 136350
rect 565274 136294 565342 136350
rect 565398 136294 565494 136350
rect 564874 136226 565494 136294
rect 564874 136170 564970 136226
rect 565026 136170 565094 136226
rect 565150 136170 565218 136226
rect 565274 136170 565342 136226
rect 565398 136170 565494 136226
rect 564874 136102 565494 136170
rect 564874 136046 564970 136102
rect 565026 136046 565094 136102
rect 565150 136046 565218 136102
rect 565274 136046 565342 136102
rect 565398 136046 565494 136102
rect 564874 135978 565494 136046
rect 564874 135922 564970 135978
rect 565026 135922 565094 135978
rect 565150 135922 565218 135978
rect 565274 135922 565342 135978
rect 565398 135922 565494 135978
rect 564874 118350 565494 135922
rect 564874 118294 564970 118350
rect 565026 118294 565094 118350
rect 565150 118294 565218 118350
rect 565274 118294 565342 118350
rect 565398 118294 565494 118350
rect 564874 118226 565494 118294
rect 564874 118170 564970 118226
rect 565026 118170 565094 118226
rect 565150 118170 565218 118226
rect 565274 118170 565342 118226
rect 565398 118170 565494 118226
rect 564874 118102 565494 118170
rect 564874 118046 564970 118102
rect 565026 118046 565094 118102
rect 565150 118046 565218 118102
rect 565274 118046 565342 118102
rect 565398 118046 565494 118102
rect 564874 117978 565494 118046
rect 564874 117922 564970 117978
rect 565026 117922 565094 117978
rect 565150 117922 565218 117978
rect 565274 117922 565342 117978
rect 565398 117922 565494 117978
rect 564874 100350 565494 117922
rect 564874 100294 564970 100350
rect 565026 100294 565094 100350
rect 565150 100294 565218 100350
rect 565274 100294 565342 100350
rect 565398 100294 565494 100350
rect 564874 100226 565494 100294
rect 564874 100170 564970 100226
rect 565026 100170 565094 100226
rect 565150 100170 565218 100226
rect 565274 100170 565342 100226
rect 565398 100170 565494 100226
rect 564874 100102 565494 100170
rect 564874 100046 564970 100102
rect 565026 100046 565094 100102
rect 565150 100046 565218 100102
rect 565274 100046 565342 100102
rect 565398 100046 565494 100102
rect 564874 99978 565494 100046
rect 564874 99922 564970 99978
rect 565026 99922 565094 99978
rect 565150 99922 565218 99978
rect 565274 99922 565342 99978
rect 565398 99922 565494 99978
rect 564874 82350 565494 99922
rect 564874 82294 564970 82350
rect 565026 82294 565094 82350
rect 565150 82294 565218 82350
rect 565274 82294 565342 82350
rect 565398 82294 565494 82350
rect 564874 82226 565494 82294
rect 564874 82170 564970 82226
rect 565026 82170 565094 82226
rect 565150 82170 565218 82226
rect 565274 82170 565342 82226
rect 565398 82170 565494 82226
rect 564874 82102 565494 82170
rect 564874 82046 564970 82102
rect 565026 82046 565094 82102
rect 565150 82046 565218 82102
rect 565274 82046 565342 82102
rect 565398 82046 565494 82102
rect 564874 81978 565494 82046
rect 564874 81922 564970 81978
rect 565026 81922 565094 81978
rect 565150 81922 565218 81978
rect 565274 81922 565342 81978
rect 565398 81922 565494 81978
rect 564874 64350 565494 81922
rect 564874 64294 564970 64350
rect 565026 64294 565094 64350
rect 565150 64294 565218 64350
rect 565274 64294 565342 64350
rect 565398 64294 565494 64350
rect 564874 64226 565494 64294
rect 564874 64170 564970 64226
rect 565026 64170 565094 64226
rect 565150 64170 565218 64226
rect 565274 64170 565342 64226
rect 565398 64170 565494 64226
rect 564874 64102 565494 64170
rect 564874 64046 564970 64102
rect 565026 64046 565094 64102
rect 565150 64046 565218 64102
rect 565274 64046 565342 64102
rect 565398 64046 565494 64102
rect 564874 63978 565494 64046
rect 564874 63922 564970 63978
rect 565026 63922 565094 63978
rect 565150 63922 565218 63978
rect 565274 63922 565342 63978
rect 565398 63922 565494 63978
rect 564874 46350 565494 63922
rect 564874 46294 564970 46350
rect 565026 46294 565094 46350
rect 565150 46294 565218 46350
rect 565274 46294 565342 46350
rect 565398 46294 565494 46350
rect 564874 46226 565494 46294
rect 564874 46170 564970 46226
rect 565026 46170 565094 46226
rect 565150 46170 565218 46226
rect 565274 46170 565342 46226
rect 565398 46170 565494 46226
rect 564874 46102 565494 46170
rect 564874 46046 564970 46102
rect 565026 46046 565094 46102
rect 565150 46046 565218 46102
rect 565274 46046 565342 46102
rect 565398 46046 565494 46102
rect 564874 45978 565494 46046
rect 564874 45922 564970 45978
rect 565026 45922 565094 45978
rect 565150 45922 565218 45978
rect 565274 45922 565342 45978
rect 565398 45922 565494 45978
rect 564874 28350 565494 45922
rect 564874 28294 564970 28350
rect 565026 28294 565094 28350
rect 565150 28294 565218 28350
rect 565274 28294 565342 28350
rect 565398 28294 565494 28350
rect 564874 28226 565494 28294
rect 564874 28170 564970 28226
rect 565026 28170 565094 28226
rect 565150 28170 565218 28226
rect 565274 28170 565342 28226
rect 565398 28170 565494 28226
rect 564874 28102 565494 28170
rect 564874 28046 564970 28102
rect 565026 28046 565094 28102
rect 565150 28046 565218 28102
rect 565274 28046 565342 28102
rect 565398 28046 565494 28102
rect 564874 27978 565494 28046
rect 564874 27922 564970 27978
rect 565026 27922 565094 27978
rect 565150 27922 565218 27978
rect 565274 27922 565342 27978
rect 565398 27922 565494 27978
rect 564874 10350 565494 27922
rect 564874 10294 564970 10350
rect 565026 10294 565094 10350
rect 565150 10294 565218 10350
rect 565274 10294 565342 10350
rect 565398 10294 565494 10350
rect 564874 10226 565494 10294
rect 564874 10170 564970 10226
rect 565026 10170 565094 10226
rect 565150 10170 565218 10226
rect 565274 10170 565342 10226
rect 565398 10170 565494 10226
rect 564874 10102 565494 10170
rect 564874 10046 564970 10102
rect 565026 10046 565094 10102
rect 565150 10046 565218 10102
rect 565274 10046 565342 10102
rect 565398 10046 565494 10102
rect 564874 9978 565494 10046
rect 564874 9922 564970 9978
rect 565026 9922 565094 9978
rect 565150 9922 565218 9978
rect 565274 9922 565342 9978
rect 565398 9922 565494 9978
rect 564874 -1120 565494 9922
rect 564874 -1176 564970 -1120
rect 565026 -1176 565094 -1120
rect 565150 -1176 565218 -1120
rect 565274 -1176 565342 -1120
rect 565398 -1176 565494 -1120
rect 564874 -1244 565494 -1176
rect 564874 -1300 564970 -1244
rect 565026 -1300 565094 -1244
rect 565150 -1300 565218 -1244
rect 565274 -1300 565342 -1244
rect 565398 -1300 565494 -1244
rect 564874 -1368 565494 -1300
rect 564874 -1424 564970 -1368
rect 565026 -1424 565094 -1368
rect 565150 -1424 565218 -1368
rect 565274 -1424 565342 -1368
rect 565398 -1424 565494 -1368
rect 564874 -1492 565494 -1424
rect 564874 -1548 564970 -1492
rect 565026 -1548 565094 -1492
rect 565150 -1548 565218 -1492
rect 565274 -1548 565342 -1492
rect 565398 -1548 565494 -1492
rect 564874 -1644 565494 -1548
rect 579154 597212 579774 598268
rect 579154 597156 579250 597212
rect 579306 597156 579374 597212
rect 579430 597156 579498 597212
rect 579554 597156 579622 597212
rect 579678 597156 579774 597212
rect 579154 597088 579774 597156
rect 579154 597032 579250 597088
rect 579306 597032 579374 597088
rect 579430 597032 579498 597088
rect 579554 597032 579622 597088
rect 579678 597032 579774 597088
rect 579154 596964 579774 597032
rect 579154 596908 579250 596964
rect 579306 596908 579374 596964
rect 579430 596908 579498 596964
rect 579554 596908 579622 596964
rect 579678 596908 579774 596964
rect 579154 596840 579774 596908
rect 579154 596784 579250 596840
rect 579306 596784 579374 596840
rect 579430 596784 579498 596840
rect 579554 596784 579622 596840
rect 579678 596784 579774 596840
rect 579154 580350 579774 596784
rect 579154 580294 579250 580350
rect 579306 580294 579374 580350
rect 579430 580294 579498 580350
rect 579554 580294 579622 580350
rect 579678 580294 579774 580350
rect 579154 580226 579774 580294
rect 579154 580170 579250 580226
rect 579306 580170 579374 580226
rect 579430 580170 579498 580226
rect 579554 580170 579622 580226
rect 579678 580170 579774 580226
rect 579154 580102 579774 580170
rect 579154 580046 579250 580102
rect 579306 580046 579374 580102
rect 579430 580046 579498 580102
rect 579554 580046 579622 580102
rect 579678 580046 579774 580102
rect 579154 579978 579774 580046
rect 579154 579922 579250 579978
rect 579306 579922 579374 579978
rect 579430 579922 579498 579978
rect 579554 579922 579622 579978
rect 579678 579922 579774 579978
rect 579154 562350 579774 579922
rect 579154 562294 579250 562350
rect 579306 562294 579374 562350
rect 579430 562294 579498 562350
rect 579554 562294 579622 562350
rect 579678 562294 579774 562350
rect 579154 562226 579774 562294
rect 579154 562170 579250 562226
rect 579306 562170 579374 562226
rect 579430 562170 579498 562226
rect 579554 562170 579622 562226
rect 579678 562170 579774 562226
rect 579154 562102 579774 562170
rect 579154 562046 579250 562102
rect 579306 562046 579374 562102
rect 579430 562046 579498 562102
rect 579554 562046 579622 562102
rect 579678 562046 579774 562102
rect 579154 561978 579774 562046
rect 579154 561922 579250 561978
rect 579306 561922 579374 561978
rect 579430 561922 579498 561978
rect 579554 561922 579622 561978
rect 579678 561922 579774 561978
rect 579154 544350 579774 561922
rect 579154 544294 579250 544350
rect 579306 544294 579374 544350
rect 579430 544294 579498 544350
rect 579554 544294 579622 544350
rect 579678 544294 579774 544350
rect 579154 544226 579774 544294
rect 579154 544170 579250 544226
rect 579306 544170 579374 544226
rect 579430 544170 579498 544226
rect 579554 544170 579622 544226
rect 579678 544170 579774 544226
rect 579154 544102 579774 544170
rect 579154 544046 579250 544102
rect 579306 544046 579374 544102
rect 579430 544046 579498 544102
rect 579554 544046 579622 544102
rect 579678 544046 579774 544102
rect 579154 543978 579774 544046
rect 579154 543922 579250 543978
rect 579306 543922 579374 543978
rect 579430 543922 579498 543978
rect 579554 543922 579622 543978
rect 579678 543922 579774 543978
rect 579154 526350 579774 543922
rect 579154 526294 579250 526350
rect 579306 526294 579374 526350
rect 579430 526294 579498 526350
rect 579554 526294 579622 526350
rect 579678 526294 579774 526350
rect 579154 526226 579774 526294
rect 579154 526170 579250 526226
rect 579306 526170 579374 526226
rect 579430 526170 579498 526226
rect 579554 526170 579622 526226
rect 579678 526170 579774 526226
rect 579154 526102 579774 526170
rect 579154 526046 579250 526102
rect 579306 526046 579374 526102
rect 579430 526046 579498 526102
rect 579554 526046 579622 526102
rect 579678 526046 579774 526102
rect 579154 525978 579774 526046
rect 579154 525922 579250 525978
rect 579306 525922 579374 525978
rect 579430 525922 579498 525978
rect 579554 525922 579622 525978
rect 579678 525922 579774 525978
rect 579154 508350 579774 525922
rect 579154 508294 579250 508350
rect 579306 508294 579374 508350
rect 579430 508294 579498 508350
rect 579554 508294 579622 508350
rect 579678 508294 579774 508350
rect 579154 508226 579774 508294
rect 579154 508170 579250 508226
rect 579306 508170 579374 508226
rect 579430 508170 579498 508226
rect 579554 508170 579622 508226
rect 579678 508170 579774 508226
rect 579154 508102 579774 508170
rect 579154 508046 579250 508102
rect 579306 508046 579374 508102
rect 579430 508046 579498 508102
rect 579554 508046 579622 508102
rect 579678 508046 579774 508102
rect 579154 507978 579774 508046
rect 579154 507922 579250 507978
rect 579306 507922 579374 507978
rect 579430 507922 579498 507978
rect 579554 507922 579622 507978
rect 579678 507922 579774 507978
rect 579154 490350 579774 507922
rect 579154 490294 579250 490350
rect 579306 490294 579374 490350
rect 579430 490294 579498 490350
rect 579554 490294 579622 490350
rect 579678 490294 579774 490350
rect 579154 490226 579774 490294
rect 579154 490170 579250 490226
rect 579306 490170 579374 490226
rect 579430 490170 579498 490226
rect 579554 490170 579622 490226
rect 579678 490170 579774 490226
rect 579154 490102 579774 490170
rect 579154 490046 579250 490102
rect 579306 490046 579374 490102
rect 579430 490046 579498 490102
rect 579554 490046 579622 490102
rect 579678 490046 579774 490102
rect 579154 489978 579774 490046
rect 579154 489922 579250 489978
rect 579306 489922 579374 489978
rect 579430 489922 579498 489978
rect 579554 489922 579622 489978
rect 579678 489922 579774 489978
rect 579154 472350 579774 489922
rect 579154 472294 579250 472350
rect 579306 472294 579374 472350
rect 579430 472294 579498 472350
rect 579554 472294 579622 472350
rect 579678 472294 579774 472350
rect 579154 472226 579774 472294
rect 579154 472170 579250 472226
rect 579306 472170 579374 472226
rect 579430 472170 579498 472226
rect 579554 472170 579622 472226
rect 579678 472170 579774 472226
rect 579154 472102 579774 472170
rect 579154 472046 579250 472102
rect 579306 472046 579374 472102
rect 579430 472046 579498 472102
rect 579554 472046 579622 472102
rect 579678 472046 579774 472102
rect 579154 471978 579774 472046
rect 579154 471922 579250 471978
rect 579306 471922 579374 471978
rect 579430 471922 579498 471978
rect 579554 471922 579622 471978
rect 579678 471922 579774 471978
rect 579154 454350 579774 471922
rect 579154 454294 579250 454350
rect 579306 454294 579374 454350
rect 579430 454294 579498 454350
rect 579554 454294 579622 454350
rect 579678 454294 579774 454350
rect 579154 454226 579774 454294
rect 579154 454170 579250 454226
rect 579306 454170 579374 454226
rect 579430 454170 579498 454226
rect 579554 454170 579622 454226
rect 579678 454170 579774 454226
rect 579154 454102 579774 454170
rect 579154 454046 579250 454102
rect 579306 454046 579374 454102
rect 579430 454046 579498 454102
rect 579554 454046 579622 454102
rect 579678 454046 579774 454102
rect 579154 453978 579774 454046
rect 579154 453922 579250 453978
rect 579306 453922 579374 453978
rect 579430 453922 579498 453978
rect 579554 453922 579622 453978
rect 579678 453922 579774 453978
rect 579154 436350 579774 453922
rect 579154 436294 579250 436350
rect 579306 436294 579374 436350
rect 579430 436294 579498 436350
rect 579554 436294 579622 436350
rect 579678 436294 579774 436350
rect 579154 436226 579774 436294
rect 579154 436170 579250 436226
rect 579306 436170 579374 436226
rect 579430 436170 579498 436226
rect 579554 436170 579622 436226
rect 579678 436170 579774 436226
rect 579154 436102 579774 436170
rect 579154 436046 579250 436102
rect 579306 436046 579374 436102
rect 579430 436046 579498 436102
rect 579554 436046 579622 436102
rect 579678 436046 579774 436102
rect 579154 435978 579774 436046
rect 579154 435922 579250 435978
rect 579306 435922 579374 435978
rect 579430 435922 579498 435978
rect 579554 435922 579622 435978
rect 579678 435922 579774 435978
rect 579154 418350 579774 435922
rect 579154 418294 579250 418350
rect 579306 418294 579374 418350
rect 579430 418294 579498 418350
rect 579554 418294 579622 418350
rect 579678 418294 579774 418350
rect 579154 418226 579774 418294
rect 579154 418170 579250 418226
rect 579306 418170 579374 418226
rect 579430 418170 579498 418226
rect 579554 418170 579622 418226
rect 579678 418170 579774 418226
rect 579154 418102 579774 418170
rect 579154 418046 579250 418102
rect 579306 418046 579374 418102
rect 579430 418046 579498 418102
rect 579554 418046 579622 418102
rect 579678 418046 579774 418102
rect 579154 417978 579774 418046
rect 579154 417922 579250 417978
rect 579306 417922 579374 417978
rect 579430 417922 579498 417978
rect 579554 417922 579622 417978
rect 579678 417922 579774 417978
rect 579154 400350 579774 417922
rect 579154 400294 579250 400350
rect 579306 400294 579374 400350
rect 579430 400294 579498 400350
rect 579554 400294 579622 400350
rect 579678 400294 579774 400350
rect 579154 400226 579774 400294
rect 579154 400170 579250 400226
rect 579306 400170 579374 400226
rect 579430 400170 579498 400226
rect 579554 400170 579622 400226
rect 579678 400170 579774 400226
rect 579154 400102 579774 400170
rect 579154 400046 579250 400102
rect 579306 400046 579374 400102
rect 579430 400046 579498 400102
rect 579554 400046 579622 400102
rect 579678 400046 579774 400102
rect 579154 399978 579774 400046
rect 579154 399922 579250 399978
rect 579306 399922 579374 399978
rect 579430 399922 579498 399978
rect 579554 399922 579622 399978
rect 579678 399922 579774 399978
rect 579154 382350 579774 399922
rect 579154 382294 579250 382350
rect 579306 382294 579374 382350
rect 579430 382294 579498 382350
rect 579554 382294 579622 382350
rect 579678 382294 579774 382350
rect 579154 382226 579774 382294
rect 579154 382170 579250 382226
rect 579306 382170 579374 382226
rect 579430 382170 579498 382226
rect 579554 382170 579622 382226
rect 579678 382170 579774 382226
rect 579154 382102 579774 382170
rect 579154 382046 579250 382102
rect 579306 382046 579374 382102
rect 579430 382046 579498 382102
rect 579554 382046 579622 382102
rect 579678 382046 579774 382102
rect 579154 381978 579774 382046
rect 579154 381922 579250 381978
rect 579306 381922 579374 381978
rect 579430 381922 579498 381978
rect 579554 381922 579622 381978
rect 579678 381922 579774 381978
rect 579154 364350 579774 381922
rect 579154 364294 579250 364350
rect 579306 364294 579374 364350
rect 579430 364294 579498 364350
rect 579554 364294 579622 364350
rect 579678 364294 579774 364350
rect 579154 364226 579774 364294
rect 579154 364170 579250 364226
rect 579306 364170 579374 364226
rect 579430 364170 579498 364226
rect 579554 364170 579622 364226
rect 579678 364170 579774 364226
rect 579154 364102 579774 364170
rect 579154 364046 579250 364102
rect 579306 364046 579374 364102
rect 579430 364046 579498 364102
rect 579554 364046 579622 364102
rect 579678 364046 579774 364102
rect 579154 363978 579774 364046
rect 579154 363922 579250 363978
rect 579306 363922 579374 363978
rect 579430 363922 579498 363978
rect 579554 363922 579622 363978
rect 579678 363922 579774 363978
rect 579154 346350 579774 363922
rect 579154 346294 579250 346350
rect 579306 346294 579374 346350
rect 579430 346294 579498 346350
rect 579554 346294 579622 346350
rect 579678 346294 579774 346350
rect 579154 346226 579774 346294
rect 579154 346170 579250 346226
rect 579306 346170 579374 346226
rect 579430 346170 579498 346226
rect 579554 346170 579622 346226
rect 579678 346170 579774 346226
rect 579154 346102 579774 346170
rect 579154 346046 579250 346102
rect 579306 346046 579374 346102
rect 579430 346046 579498 346102
rect 579554 346046 579622 346102
rect 579678 346046 579774 346102
rect 579154 345978 579774 346046
rect 579154 345922 579250 345978
rect 579306 345922 579374 345978
rect 579430 345922 579498 345978
rect 579554 345922 579622 345978
rect 579678 345922 579774 345978
rect 579154 328350 579774 345922
rect 579154 328294 579250 328350
rect 579306 328294 579374 328350
rect 579430 328294 579498 328350
rect 579554 328294 579622 328350
rect 579678 328294 579774 328350
rect 579154 328226 579774 328294
rect 579154 328170 579250 328226
rect 579306 328170 579374 328226
rect 579430 328170 579498 328226
rect 579554 328170 579622 328226
rect 579678 328170 579774 328226
rect 579154 328102 579774 328170
rect 579154 328046 579250 328102
rect 579306 328046 579374 328102
rect 579430 328046 579498 328102
rect 579554 328046 579622 328102
rect 579678 328046 579774 328102
rect 579154 327978 579774 328046
rect 579154 327922 579250 327978
rect 579306 327922 579374 327978
rect 579430 327922 579498 327978
rect 579554 327922 579622 327978
rect 579678 327922 579774 327978
rect 579154 310350 579774 327922
rect 579154 310294 579250 310350
rect 579306 310294 579374 310350
rect 579430 310294 579498 310350
rect 579554 310294 579622 310350
rect 579678 310294 579774 310350
rect 579154 310226 579774 310294
rect 579154 310170 579250 310226
rect 579306 310170 579374 310226
rect 579430 310170 579498 310226
rect 579554 310170 579622 310226
rect 579678 310170 579774 310226
rect 579154 310102 579774 310170
rect 579154 310046 579250 310102
rect 579306 310046 579374 310102
rect 579430 310046 579498 310102
rect 579554 310046 579622 310102
rect 579678 310046 579774 310102
rect 579154 309978 579774 310046
rect 579154 309922 579250 309978
rect 579306 309922 579374 309978
rect 579430 309922 579498 309978
rect 579554 309922 579622 309978
rect 579678 309922 579774 309978
rect 579154 292350 579774 309922
rect 579154 292294 579250 292350
rect 579306 292294 579374 292350
rect 579430 292294 579498 292350
rect 579554 292294 579622 292350
rect 579678 292294 579774 292350
rect 579154 292226 579774 292294
rect 579154 292170 579250 292226
rect 579306 292170 579374 292226
rect 579430 292170 579498 292226
rect 579554 292170 579622 292226
rect 579678 292170 579774 292226
rect 579154 292102 579774 292170
rect 579154 292046 579250 292102
rect 579306 292046 579374 292102
rect 579430 292046 579498 292102
rect 579554 292046 579622 292102
rect 579678 292046 579774 292102
rect 579154 291978 579774 292046
rect 579154 291922 579250 291978
rect 579306 291922 579374 291978
rect 579430 291922 579498 291978
rect 579554 291922 579622 291978
rect 579678 291922 579774 291978
rect 579154 274350 579774 291922
rect 579154 274294 579250 274350
rect 579306 274294 579374 274350
rect 579430 274294 579498 274350
rect 579554 274294 579622 274350
rect 579678 274294 579774 274350
rect 579154 274226 579774 274294
rect 579154 274170 579250 274226
rect 579306 274170 579374 274226
rect 579430 274170 579498 274226
rect 579554 274170 579622 274226
rect 579678 274170 579774 274226
rect 579154 274102 579774 274170
rect 579154 274046 579250 274102
rect 579306 274046 579374 274102
rect 579430 274046 579498 274102
rect 579554 274046 579622 274102
rect 579678 274046 579774 274102
rect 579154 273978 579774 274046
rect 579154 273922 579250 273978
rect 579306 273922 579374 273978
rect 579430 273922 579498 273978
rect 579554 273922 579622 273978
rect 579678 273922 579774 273978
rect 579154 256350 579774 273922
rect 579154 256294 579250 256350
rect 579306 256294 579374 256350
rect 579430 256294 579498 256350
rect 579554 256294 579622 256350
rect 579678 256294 579774 256350
rect 579154 256226 579774 256294
rect 579154 256170 579250 256226
rect 579306 256170 579374 256226
rect 579430 256170 579498 256226
rect 579554 256170 579622 256226
rect 579678 256170 579774 256226
rect 579154 256102 579774 256170
rect 579154 256046 579250 256102
rect 579306 256046 579374 256102
rect 579430 256046 579498 256102
rect 579554 256046 579622 256102
rect 579678 256046 579774 256102
rect 579154 255978 579774 256046
rect 579154 255922 579250 255978
rect 579306 255922 579374 255978
rect 579430 255922 579498 255978
rect 579554 255922 579622 255978
rect 579678 255922 579774 255978
rect 579154 238350 579774 255922
rect 579154 238294 579250 238350
rect 579306 238294 579374 238350
rect 579430 238294 579498 238350
rect 579554 238294 579622 238350
rect 579678 238294 579774 238350
rect 579154 238226 579774 238294
rect 579154 238170 579250 238226
rect 579306 238170 579374 238226
rect 579430 238170 579498 238226
rect 579554 238170 579622 238226
rect 579678 238170 579774 238226
rect 579154 238102 579774 238170
rect 579154 238046 579250 238102
rect 579306 238046 579374 238102
rect 579430 238046 579498 238102
rect 579554 238046 579622 238102
rect 579678 238046 579774 238102
rect 579154 237978 579774 238046
rect 579154 237922 579250 237978
rect 579306 237922 579374 237978
rect 579430 237922 579498 237978
rect 579554 237922 579622 237978
rect 579678 237922 579774 237978
rect 579154 220350 579774 237922
rect 579154 220294 579250 220350
rect 579306 220294 579374 220350
rect 579430 220294 579498 220350
rect 579554 220294 579622 220350
rect 579678 220294 579774 220350
rect 579154 220226 579774 220294
rect 579154 220170 579250 220226
rect 579306 220170 579374 220226
rect 579430 220170 579498 220226
rect 579554 220170 579622 220226
rect 579678 220170 579774 220226
rect 579154 220102 579774 220170
rect 579154 220046 579250 220102
rect 579306 220046 579374 220102
rect 579430 220046 579498 220102
rect 579554 220046 579622 220102
rect 579678 220046 579774 220102
rect 579154 219978 579774 220046
rect 579154 219922 579250 219978
rect 579306 219922 579374 219978
rect 579430 219922 579498 219978
rect 579554 219922 579622 219978
rect 579678 219922 579774 219978
rect 579154 202350 579774 219922
rect 579154 202294 579250 202350
rect 579306 202294 579374 202350
rect 579430 202294 579498 202350
rect 579554 202294 579622 202350
rect 579678 202294 579774 202350
rect 579154 202226 579774 202294
rect 579154 202170 579250 202226
rect 579306 202170 579374 202226
rect 579430 202170 579498 202226
rect 579554 202170 579622 202226
rect 579678 202170 579774 202226
rect 579154 202102 579774 202170
rect 579154 202046 579250 202102
rect 579306 202046 579374 202102
rect 579430 202046 579498 202102
rect 579554 202046 579622 202102
rect 579678 202046 579774 202102
rect 579154 201978 579774 202046
rect 579154 201922 579250 201978
rect 579306 201922 579374 201978
rect 579430 201922 579498 201978
rect 579554 201922 579622 201978
rect 579678 201922 579774 201978
rect 579154 184350 579774 201922
rect 579154 184294 579250 184350
rect 579306 184294 579374 184350
rect 579430 184294 579498 184350
rect 579554 184294 579622 184350
rect 579678 184294 579774 184350
rect 579154 184226 579774 184294
rect 579154 184170 579250 184226
rect 579306 184170 579374 184226
rect 579430 184170 579498 184226
rect 579554 184170 579622 184226
rect 579678 184170 579774 184226
rect 579154 184102 579774 184170
rect 579154 184046 579250 184102
rect 579306 184046 579374 184102
rect 579430 184046 579498 184102
rect 579554 184046 579622 184102
rect 579678 184046 579774 184102
rect 579154 183978 579774 184046
rect 579154 183922 579250 183978
rect 579306 183922 579374 183978
rect 579430 183922 579498 183978
rect 579554 183922 579622 183978
rect 579678 183922 579774 183978
rect 579154 166350 579774 183922
rect 579154 166294 579250 166350
rect 579306 166294 579374 166350
rect 579430 166294 579498 166350
rect 579554 166294 579622 166350
rect 579678 166294 579774 166350
rect 579154 166226 579774 166294
rect 579154 166170 579250 166226
rect 579306 166170 579374 166226
rect 579430 166170 579498 166226
rect 579554 166170 579622 166226
rect 579678 166170 579774 166226
rect 579154 166102 579774 166170
rect 579154 166046 579250 166102
rect 579306 166046 579374 166102
rect 579430 166046 579498 166102
rect 579554 166046 579622 166102
rect 579678 166046 579774 166102
rect 579154 165978 579774 166046
rect 579154 165922 579250 165978
rect 579306 165922 579374 165978
rect 579430 165922 579498 165978
rect 579554 165922 579622 165978
rect 579678 165922 579774 165978
rect 579154 148350 579774 165922
rect 579154 148294 579250 148350
rect 579306 148294 579374 148350
rect 579430 148294 579498 148350
rect 579554 148294 579622 148350
rect 579678 148294 579774 148350
rect 579154 148226 579774 148294
rect 579154 148170 579250 148226
rect 579306 148170 579374 148226
rect 579430 148170 579498 148226
rect 579554 148170 579622 148226
rect 579678 148170 579774 148226
rect 579154 148102 579774 148170
rect 579154 148046 579250 148102
rect 579306 148046 579374 148102
rect 579430 148046 579498 148102
rect 579554 148046 579622 148102
rect 579678 148046 579774 148102
rect 579154 147978 579774 148046
rect 579154 147922 579250 147978
rect 579306 147922 579374 147978
rect 579430 147922 579498 147978
rect 579554 147922 579622 147978
rect 579678 147922 579774 147978
rect 579154 130350 579774 147922
rect 579154 130294 579250 130350
rect 579306 130294 579374 130350
rect 579430 130294 579498 130350
rect 579554 130294 579622 130350
rect 579678 130294 579774 130350
rect 579154 130226 579774 130294
rect 579154 130170 579250 130226
rect 579306 130170 579374 130226
rect 579430 130170 579498 130226
rect 579554 130170 579622 130226
rect 579678 130170 579774 130226
rect 579154 130102 579774 130170
rect 579154 130046 579250 130102
rect 579306 130046 579374 130102
rect 579430 130046 579498 130102
rect 579554 130046 579622 130102
rect 579678 130046 579774 130102
rect 579154 129978 579774 130046
rect 579154 129922 579250 129978
rect 579306 129922 579374 129978
rect 579430 129922 579498 129978
rect 579554 129922 579622 129978
rect 579678 129922 579774 129978
rect 579154 112350 579774 129922
rect 579154 112294 579250 112350
rect 579306 112294 579374 112350
rect 579430 112294 579498 112350
rect 579554 112294 579622 112350
rect 579678 112294 579774 112350
rect 579154 112226 579774 112294
rect 579154 112170 579250 112226
rect 579306 112170 579374 112226
rect 579430 112170 579498 112226
rect 579554 112170 579622 112226
rect 579678 112170 579774 112226
rect 579154 112102 579774 112170
rect 579154 112046 579250 112102
rect 579306 112046 579374 112102
rect 579430 112046 579498 112102
rect 579554 112046 579622 112102
rect 579678 112046 579774 112102
rect 579154 111978 579774 112046
rect 579154 111922 579250 111978
rect 579306 111922 579374 111978
rect 579430 111922 579498 111978
rect 579554 111922 579622 111978
rect 579678 111922 579774 111978
rect 579154 94350 579774 111922
rect 579154 94294 579250 94350
rect 579306 94294 579374 94350
rect 579430 94294 579498 94350
rect 579554 94294 579622 94350
rect 579678 94294 579774 94350
rect 579154 94226 579774 94294
rect 579154 94170 579250 94226
rect 579306 94170 579374 94226
rect 579430 94170 579498 94226
rect 579554 94170 579622 94226
rect 579678 94170 579774 94226
rect 579154 94102 579774 94170
rect 579154 94046 579250 94102
rect 579306 94046 579374 94102
rect 579430 94046 579498 94102
rect 579554 94046 579622 94102
rect 579678 94046 579774 94102
rect 579154 93978 579774 94046
rect 579154 93922 579250 93978
rect 579306 93922 579374 93978
rect 579430 93922 579498 93978
rect 579554 93922 579622 93978
rect 579678 93922 579774 93978
rect 579154 76350 579774 93922
rect 579154 76294 579250 76350
rect 579306 76294 579374 76350
rect 579430 76294 579498 76350
rect 579554 76294 579622 76350
rect 579678 76294 579774 76350
rect 579154 76226 579774 76294
rect 579154 76170 579250 76226
rect 579306 76170 579374 76226
rect 579430 76170 579498 76226
rect 579554 76170 579622 76226
rect 579678 76170 579774 76226
rect 579154 76102 579774 76170
rect 579154 76046 579250 76102
rect 579306 76046 579374 76102
rect 579430 76046 579498 76102
rect 579554 76046 579622 76102
rect 579678 76046 579774 76102
rect 579154 75978 579774 76046
rect 579154 75922 579250 75978
rect 579306 75922 579374 75978
rect 579430 75922 579498 75978
rect 579554 75922 579622 75978
rect 579678 75922 579774 75978
rect 579154 58350 579774 75922
rect 579154 58294 579250 58350
rect 579306 58294 579374 58350
rect 579430 58294 579498 58350
rect 579554 58294 579622 58350
rect 579678 58294 579774 58350
rect 579154 58226 579774 58294
rect 579154 58170 579250 58226
rect 579306 58170 579374 58226
rect 579430 58170 579498 58226
rect 579554 58170 579622 58226
rect 579678 58170 579774 58226
rect 579154 58102 579774 58170
rect 579154 58046 579250 58102
rect 579306 58046 579374 58102
rect 579430 58046 579498 58102
rect 579554 58046 579622 58102
rect 579678 58046 579774 58102
rect 579154 57978 579774 58046
rect 579154 57922 579250 57978
rect 579306 57922 579374 57978
rect 579430 57922 579498 57978
rect 579554 57922 579622 57978
rect 579678 57922 579774 57978
rect 579154 40350 579774 57922
rect 579154 40294 579250 40350
rect 579306 40294 579374 40350
rect 579430 40294 579498 40350
rect 579554 40294 579622 40350
rect 579678 40294 579774 40350
rect 579154 40226 579774 40294
rect 579154 40170 579250 40226
rect 579306 40170 579374 40226
rect 579430 40170 579498 40226
rect 579554 40170 579622 40226
rect 579678 40170 579774 40226
rect 579154 40102 579774 40170
rect 579154 40046 579250 40102
rect 579306 40046 579374 40102
rect 579430 40046 579498 40102
rect 579554 40046 579622 40102
rect 579678 40046 579774 40102
rect 579154 39978 579774 40046
rect 579154 39922 579250 39978
rect 579306 39922 579374 39978
rect 579430 39922 579498 39978
rect 579554 39922 579622 39978
rect 579678 39922 579774 39978
rect 579154 22350 579774 39922
rect 579154 22294 579250 22350
rect 579306 22294 579374 22350
rect 579430 22294 579498 22350
rect 579554 22294 579622 22350
rect 579678 22294 579774 22350
rect 579154 22226 579774 22294
rect 579154 22170 579250 22226
rect 579306 22170 579374 22226
rect 579430 22170 579498 22226
rect 579554 22170 579622 22226
rect 579678 22170 579774 22226
rect 579154 22102 579774 22170
rect 579154 22046 579250 22102
rect 579306 22046 579374 22102
rect 579430 22046 579498 22102
rect 579554 22046 579622 22102
rect 579678 22046 579774 22102
rect 579154 21978 579774 22046
rect 579154 21922 579250 21978
rect 579306 21922 579374 21978
rect 579430 21922 579498 21978
rect 579554 21922 579622 21978
rect 579678 21922 579774 21978
rect 579154 4350 579774 21922
rect 579154 4294 579250 4350
rect 579306 4294 579374 4350
rect 579430 4294 579498 4350
rect 579554 4294 579622 4350
rect 579678 4294 579774 4350
rect 579154 4226 579774 4294
rect 579154 4170 579250 4226
rect 579306 4170 579374 4226
rect 579430 4170 579498 4226
rect 579554 4170 579622 4226
rect 579678 4170 579774 4226
rect 579154 4102 579774 4170
rect 579154 4046 579250 4102
rect 579306 4046 579374 4102
rect 579430 4046 579498 4102
rect 579554 4046 579622 4102
rect 579678 4046 579774 4102
rect 579154 3978 579774 4046
rect 579154 3922 579250 3978
rect 579306 3922 579374 3978
rect 579430 3922 579498 3978
rect 579554 3922 579622 3978
rect 579678 3922 579774 3978
rect 579154 -160 579774 3922
rect 579154 -216 579250 -160
rect 579306 -216 579374 -160
rect 579430 -216 579498 -160
rect 579554 -216 579622 -160
rect 579678 -216 579774 -160
rect 579154 -284 579774 -216
rect 579154 -340 579250 -284
rect 579306 -340 579374 -284
rect 579430 -340 579498 -284
rect 579554 -340 579622 -284
rect 579678 -340 579774 -284
rect 579154 -408 579774 -340
rect 579154 -464 579250 -408
rect 579306 -464 579374 -408
rect 579430 -464 579498 -408
rect 579554 -464 579622 -408
rect 579678 -464 579774 -408
rect 579154 -532 579774 -464
rect 579154 -588 579250 -532
rect 579306 -588 579374 -532
rect 579430 -588 579498 -532
rect 579554 -588 579622 -532
rect 579678 -588 579774 -532
rect 579154 -1644 579774 -588
rect 582874 598172 583494 598268
rect 582874 598116 582970 598172
rect 583026 598116 583094 598172
rect 583150 598116 583218 598172
rect 583274 598116 583342 598172
rect 583398 598116 583494 598172
rect 582874 598048 583494 598116
rect 582874 597992 582970 598048
rect 583026 597992 583094 598048
rect 583150 597992 583218 598048
rect 583274 597992 583342 598048
rect 583398 597992 583494 598048
rect 582874 597924 583494 597992
rect 582874 597868 582970 597924
rect 583026 597868 583094 597924
rect 583150 597868 583218 597924
rect 583274 597868 583342 597924
rect 583398 597868 583494 597924
rect 582874 597800 583494 597868
rect 582874 597744 582970 597800
rect 583026 597744 583094 597800
rect 583150 597744 583218 597800
rect 583274 597744 583342 597800
rect 583398 597744 583494 597800
rect 582874 586350 583494 597744
rect 597360 598172 597980 598268
rect 597360 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect 597360 598048 597980 598116
rect 597360 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect 597360 597924 597980 597992
rect 597360 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect 597360 597800 597980 597868
rect 597360 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect 582874 586294 582970 586350
rect 583026 586294 583094 586350
rect 583150 586294 583218 586350
rect 583274 586294 583342 586350
rect 583398 586294 583494 586350
rect 582874 586226 583494 586294
rect 582874 586170 582970 586226
rect 583026 586170 583094 586226
rect 583150 586170 583218 586226
rect 583274 586170 583342 586226
rect 583398 586170 583494 586226
rect 582874 586102 583494 586170
rect 582874 586046 582970 586102
rect 583026 586046 583094 586102
rect 583150 586046 583218 586102
rect 583274 586046 583342 586102
rect 583398 586046 583494 586102
rect 582874 585978 583494 586046
rect 582874 585922 582970 585978
rect 583026 585922 583094 585978
rect 583150 585922 583218 585978
rect 583274 585922 583342 585978
rect 583398 585922 583494 585978
rect 582874 568350 583494 585922
rect 582874 568294 582970 568350
rect 583026 568294 583094 568350
rect 583150 568294 583218 568350
rect 583274 568294 583342 568350
rect 583398 568294 583494 568350
rect 582874 568226 583494 568294
rect 582874 568170 582970 568226
rect 583026 568170 583094 568226
rect 583150 568170 583218 568226
rect 583274 568170 583342 568226
rect 583398 568170 583494 568226
rect 582874 568102 583494 568170
rect 582874 568046 582970 568102
rect 583026 568046 583094 568102
rect 583150 568046 583218 568102
rect 583274 568046 583342 568102
rect 583398 568046 583494 568102
rect 582874 567978 583494 568046
rect 582874 567922 582970 567978
rect 583026 567922 583094 567978
rect 583150 567922 583218 567978
rect 583274 567922 583342 567978
rect 583398 567922 583494 567978
rect 582874 550350 583494 567922
rect 582874 550294 582970 550350
rect 583026 550294 583094 550350
rect 583150 550294 583218 550350
rect 583274 550294 583342 550350
rect 583398 550294 583494 550350
rect 582874 550226 583494 550294
rect 582874 550170 582970 550226
rect 583026 550170 583094 550226
rect 583150 550170 583218 550226
rect 583274 550170 583342 550226
rect 583398 550170 583494 550226
rect 582874 550102 583494 550170
rect 582874 550046 582970 550102
rect 583026 550046 583094 550102
rect 583150 550046 583218 550102
rect 583274 550046 583342 550102
rect 583398 550046 583494 550102
rect 582874 549978 583494 550046
rect 582874 549922 582970 549978
rect 583026 549922 583094 549978
rect 583150 549922 583218 549978
rect 583274 549922 583342 549978
rect 583398 549922 583494 549978
rect 582874 532350 583494 549922
rect 582874 532294 582970 532350
rect 583026 532294 583094 532350
rect 583150 532294 583218 532350
rect 583274 532294 583342 532350
rect 583398 532294 583494 532350
rect 582874 532226 583494 532294
rect 582874 532170 582970 532226
rect 583026 532170 583094 532226
rect 583150 532170 583218 532226
rect 583274 532170 583342 532226
rect 583398 532170 583494 532226
rect 582874 532102 583494 532170
rect 582874 532046 582970 532102
rect 583026 532046 583094 532102
rect 583150 532046 583218 532102
rect 583274 532046 583342 532102
rect 583398 532046 583494 532102
rect 582874 531978 583494 532046
rect 582874 531922 582970 531978
rect 583026 531922 583094 531978
rect 583150 531922 583218 531978
rect 583274 531922 583342 531978
rect 583398 531922 583494 531978
rect 582874 514350 583494 531922
rect 582874 514294 582970 514350
rect 583026 514294 583094 514350
rect 583150 514294 583218 514350
rect 583274 514294 583342 514350
rect 583398 514294 583494 514350
rect 582874 514226 583494 514294
rect 582874 514170 582970 514226
rect 583026 514170 583094 514226
rect 583150 514170 583218 514226
rect 583274 514170 583342 514226
rect 583398 514170 583494 514226
rect 582874 514102 583494 514170
rect 582874 514046 582970 514102
rect 583026 514046 583094 514102
rect 583150 514046 583218 514102
rect 583274 514046 583342 514102
rect 583398 514046 583494 514102
rect 582874 513978 583494 514046
rect 582874 513922 582970 513978
rect 583026 513922 583094 513978
rect 583150 513922 583218 513978
rect 583274 513922 583342 513978
rect 583398 513922 583494 513978
rect 582874 496350 583494 513922
rect 582874 496294 582970 496350
rect 583026 496294 583094 496350
rect 583150 496294 583218 496350
rect 583274 496294 583342 496350
rect 583398 496294 583494 496350
rect 582874 496226 583494 496294
rect 582874 496170 582970 496226
rect 583026 496170 583094 496226
rect 583150 496170 583218 496226
rect 583274 496170 583342 496226
rect 583398 496170 583494 496226
rect 582874 496102 583494 496170
rect 582874 496046 582970 496102
rect 583026 496046 583094 496102
rect 583150 496046 583218 496102
rect 583274 496046 583342 496102
rect 583398 496046 583494 496102
rect 582874 495978 583494 496046
rect 582874 495922 582970 495978
rect 583026 495922 583094 495978
rect 583150 495922 583218 495978
rect 583274 495922 583342 495978
rect 583398 495922 583494 495978
rect 582874 478350 583494 495922
rect 582874 478294 582970 478350
rect 583026 478294 583094 478350
rect 583150 478294 583218 478350
rect 583274 478294 583342 478350
rect 583398 478294 583494 478350
rect 582874 478226 583494 478294
rect 582874 478170 582970 478226
rect 583026 478170 583094 478226
rect 583150 478170 583218 478226
rect 583274 478170 583342 478226
rect 583398 478170 583494 478226
rect 582874 478102 583494 478170
rect 582874 478046 582970 478102
rect 583026 478046 583094 478102
rect 583150 478046 583218 478102
rect 583274 478046 583342 478102
rect 583398 478046 583494 478102
rect 582874 477978 583494 478046
rect 582874 477922 582970 477978
rect 583026 477922 583094 477978
rect 583150 477922 583218 477978
rect 583274 477922 583342 477978
rect 583398 477922 583494 477978
rect 582874 460350 583494 477922
rect 582874 460294 582970 460350
rect 583026 460294 583094 460350
rect 583150 460294 583218 460350
rect 583274 460294 583342 460350
rect 583398 460294 583494 460350
rect 582874 460226 583494 460294
rect 582874 460170 582970 460226
rect 583026 460170 583094 460226
rect 583150 460170 583218 460226
rect 583274 460170 583342 460226
rect 583398 460170 583494 460226
rect 582874 460102 583494 460170
rect 582874 460046 582970 460102
rect 583026 460046 583094 460102
rect 583150 460046 583218 460102
rect 583274 460046 583342 460102
rect 583398 460046 583494 460102
rect 582874 459978 583494 460046
rect 582874 459922 582970 459978
rect 583026 459922 583094 459978
rect 583150 459922 583218 459978
rect 583274 459922 583342 459978
rect 583398 459922 583494 459978
rect 582874 442350 583494 459922
rect 582874 442294 582970 442350
rect 583026 442294 583094 442350
rect 583150 442294 583218 442350
rect 583274 442294 583342 442350
rect 583398 442294 583494 442350
rect 582874 442226 583494 442294
rect 582874 442170 582970 442226
rect 583026 442170 583094 442226
rect 583150 442170 583218 442226
rect 583274 442170 583342 442226
rect 583398 442170 583494 442226
rect 582874 442102 583494 442170
rect 582874 442046 582970 442102
rect 583026 442046 583094 442102
rect 583150 442046 583218 442102
rect 583274 442046 583342 442102
rect 583398 442046 583494 442102
rect 582874 441978 583494 442046
rect 582874 441922 582970 441978
rect 583026 441922 583094 441978
rect 583150 441922 583218 441978
rect 583274 441922 583342 441978
rect 583398 441922 583494 441978
rect 582874 424350 583494 441922
rect 582874 424294 582970 424350
rect 583026 424294 583094 424350
rect 583150 424294 583218 424350
rect 583274 424294 583342 424350
rect 583398 424294 583494 424350
rect 582874 424226 583494 424294
rect 582874 424170 582970 424226
rect 583026 424170 583094 424226
rect 583150 424170 583218 424226
rect 583274 424170 583342 424226
rect 583398 424170 583494 424226
rect 582874 424102 583494 424170
rect 582874 424046 582970 424102
rect 583026 424046 583094 424102
rect 583150 424046 583218 424102
rect 583274 424046 583342 424102
rect 583398 424046 583494 424102
rect 582874 423978 583494 424046
rect 582874 423922 582970 423978
rect 583026 423922 583094 423978
rect 583150 423922 583218 423978
rect 583274 423922 583342 423978
rect 583398 423922 583494 423978
rect 582874 406350 583494 423922
rect 582874 406294 582970 406350
rect 583026 406294 583094 406350
rect 583150 406294 583218 406350
rect 583274 406294 583342 406350
rect 583398 406294 583494 406350
rect 582874 406226 583494 406294
rect 582874 406170 582970 406226
rect 583026 406170 583094 406226
rect 583150 406170 583218 406226
rect 583274 406170 583342 406226
rect 583398 406170 583494 406226
rect 582874 406102 583494 406170
rect 582874 406046 582970 406102
rect 583026 406046 583094 406102
rect 583150 406046 583218 406102
rect 583274 406046 583342 406102
rect 583398 406046 583494 406102
rect 582874 405978 583494 406046
rect 582874 405922 582970 405978
rect 583026 405922 583094 405978
rect 583150 405922 583218 405978
rect 583274 405922 583342 405978
rect 583398 405922 583494 405978
rect 582874 388350 583494 405922
rect 582874 388294 582970 388350
rect 583026 388294 583094 388350
rect 583150 388294 583218 388350
rect 583274 388294 583342 388350
rect 583398 388294 583494 388350
rect 582874 388226 583494 388294
rect 582874 388170 582970 388226
rect 583026 388170 583094 388226
rect 583150 388170 583218 388226
rect 583274 388170 583342 388226
rect 583398 388170 583494 388226
rect 582874 388102 583494 388170
rect 582874 388046 582970 388102
rect 583026 388046 583094 388102
rect 583150 388046 583218 388102
rect 583274 388046 583342 388102
rect 583398 388046 583494 388102
rect 582874 387978 583494 388046
rect 582874 387922 582970 387978
rect 583026 387922 583094 387978
rect 583150 387922 583218 387978
rect 583274 387922 583342 387978
rect 583398 387922 583494 387978
rect 582874 370350 583494 387922
rect 582874 370294 582970 370350
rect 583026 370294 583094 370350
rect 583150 370294 583218 370350
rect 583274 370294 583342 370350
rect 583398 370294 583494 370350
rect 582874 370226 583494 370294
rect 582874 370170 582970 370226
rect 583026 370170 583094 370226
rect 583150 370170 583218 370226
rect 583274 370170 583342 370226
rect 583398 370170 583494 370226
rect 582874 370102 583494 370170
rect 582874 370046 582970 370102
rect 583026 370046 583094 370102
rect 583150 370046 583218 370102
rect 583274 370046 583342 370102
rect 583398 370046 583494 370102
rect 582874 369978 583494 370046
rect 582874 369922 582970 369978
rect 583026 369922 583094 369978
rect 583150 369922 583218 369978
rect 583274 369922 583342 369978
rect 583398 369922 583494 369978
rect 582874 352350 583494 369922
rect 582874 352294 582970 352350
rect 583026 352294 583094 352350
rect 583150 352294 583218 352350
rect 583274 352294 583342 352350
rect 583398 352294 583494 352350
rect 582874 352226 583494 352294
rect 582874 352170 582970 352226
rect 583026 352170 583094 352226
rect 583150 352170 583218 352226
rect 583274 352170 583342 352226
rect 583398 352170 583494 352226
rect 582874 352102 583494 352170
rect 582874 352046 582970 352102
rect 583026 352046 583094 352102
rect 583150 352046 583218 352102
rect 583274 352046 583342 352102
rect 583398 352046 583494 352102
rect 582874 351978 583494 352046
rect 582874 351922 582970 351978
rect 583026 351922 583094 351978
rect 583150 351922 583218 351978
rect 583274 351922 583342 351978
rect 583398 351922 583494 351978
rect 582874 334350 583494 351922
rect 582874 334294 582970 334350
rect 583026 334294 583094 334350
rect 583150 334294 583218 334350
rect 583274 334294 583342 334350
rect 583398 334294 583494 334350
rect 582874 334226 583494 334294
rect 582874 334170 582970 334226
rect 583026 334170 583094 334226
rect 583150 334170 583218 334226
rect 583274 334170 583342 334226
rect 583398 334170 583494 334226
rect 582874 334102 583494 334170
rect 582874 334046 582970 334102
rect 583026 334046 583094 334102
rect 583150 334046 583218 334102
rect 583274 334046 583342 334102
rect 583398 334046 583494 334102
rect 582874 333978 583494 334046
rect 582874 333922 582970 333978
rect 583026 333922 583094 333978
rect 583150 333922 583218 333978
rect 583274 333922 583342 333978
rect 583398 333922 583494 333978
rect 582874 316350 583494 333922
rect 582874 316294 582970 316350
rect 583026 316294 583094 316350
rect 583150 316294 583218 316350
rect 583274 316294 583342 316350
rect 583398 316294 583494 316350
rect 582874 316226 583494 316294
rect 582874 316170 582970 316226
rect 583026 316170 583094 316226
rect 583150 316170 583218 316226
rect 583274 316170 583342 316226
rect 583398 316170 583494 316226
rect 582874 316102 583494 316170
rect 582874 316046 582970 316102
rect 583026 316046 583094 316102
rect 583150 316046 583218 316102
rect 583274 316046 583342 316102
rect 583398 316046 583494 316102
rect 582874 315978 583494 316046
rect 582874 315922 582970 315978
rect 583026 315922 583094 315978
rect 583150 315922 583218 315978
rect 583274 315922 583342 315978
rect 583398 315922 583494 315978
rect 582874 298350 583494 315922
rect 582874 298294 582970 298350
rect 583026 298294 583094 298350
rect 583150 298294 583218 298350
rect 583274 298294 583342 298350
rect 583398 298294 583494 298350
rect 582874 298226 583494 298294
rect 582874 298170 582970 298226
rect 583026 298170 583094 298226
rect 583150 298170 583218 298226
rect 583274 298170 583342 298226
rect 583398 298170 583494 298226
rect 582874 298102 583494 298170
rect 582874 298046 582970 298102
rect 583026 298046 583094 298102
rect 583150 298046 583218 298102
rect 583274 298046 583342 298102
rect 583398 298046 583494 298102
rect 582874 297978 583494 298046
rect 582874 297922 582970 297978
rect 583026 297922 583094 297978
rect 583150 297922 583218 297978
rect 583274 297922 583342 297978
rect 583398 297922 583494 297978
rect 582874 280350 583494 297922
rect 582874 280294 582970 280350
rect 583026 280294 583094 280350
rect 583150 280294 583218 280350
rect 583274 280294 583342 280350
rect 583398 280294 583494 280350
rect 582874 280226 583494 280294
rect 582874 280170 582970 280226
rect 583026 280170 583094 280226
rect 583150 280170 583218 280226
rect 583274 280170 583342 280226
rect 583398 280170 583494 280226
rect 582874 280102 583494 280170
rect 582874 280046 582970 280102
rect 583026 280046 583094 280102
rect 583150 280046 583218 280102
rect 583274 280046 583342 280102
rect 583398 280046 583494 280102
rect 582874 279978 583494 280046
rect 582874 279922 582970 279978
rect 583026 279922 583094 279978
rect 583150 279922 583218 279978
rect 583274 279922 583342 279978
rect 583398 279922 583494 279978
rect 582874 262350 583494 279922
rect 582874 262294 582970 262350
rect 583026 262294 583094 262350
rect 583150 262294 583218 262350
rect 583274 262294 583342 262350
rect 583398 262294 583494 262350
rect 582874 262226 583494 262294
rect 582874 262170 582970 262226
rect 583026 262170 583094 262226
rect 583150 262170 583218 262226
rect 583274 262170 583342 262226
rect 583398 262170 583494 262226
rect 582874 262102 583494 262170
rect 582874 262046 582970 262102
rect 583026 262046 583094 262102
rect 583150 262046 583218 262102
rect 583274 262046 583342 262102
rect 583398 262046 583494 262102
rect 582874 261978 583494 262046
rect 582874 261922 582970 261978
rect 583026 261922 583094 261978
rect 583150 261922 583218 261978
rect 583274 261922 583342 261978
rect 583398 261922 583494 261978
rect 582874 244350 583494 261922
rect 582874 244294 582970 244350
rect 583026 244294 583094 244350
rect 583150 244294 583218 244350
rect 583274 244294 583342 244350
rect 583398 244294 583494 244350
rect 582874 244226 583494 244294
rect 582874 244170 582970 244226
rect 583026 244170 583094 244226
rect 583150 244170 583218 244226
rect 583274 244170 583342 244226
rect 583398 244170 583494 244226
rect 582874 244102 583494 244170
rect 582874 244046 582970 244102
rect 583026 244046 583094 244102
rect 583150 244046 583218 244102
rect 583274 244046 583342 244102
rect 583398 244046 583494 244102
rect 582874 243978 583494 244046
rect 582874 243922 582970 243978
rect 583026 243922 583094 243978
rect 583150 243922 583218 243978
rect 583274 243922 583342 243978
rect 583398 243922 583494 243978
rect 582874 226350 583494 243922
rect 582874 226294 582970 226350
rect 583026 226294 583094 226350
rect 583150 226294 583218 226350
rect 583274 226294 583342 226350
rect 583398 226294 583494 226350
rect 582874 226226 583494 226294
rect 582874 226170 582970 226226
rect 583026 226170 583094 226226
rect 583150 226170 583218 226226
rect 583274 226170 583342 226226
rect 583398 226170 583494 226226
rect 582874 226102 583494 226170
rect 582874 226046 582970 226102
rect 583026 226046 583094 226102
rect 583150 226046 583218 226102
rect 583274 226046 583342 226102
rect 583398 226046 583494 226102
rect 582874 225978 583494 226046
rect 582874 225922 582970 225978
rect 583026 225922 583094 225978
rect 583150 225922 583218 225978
rect 583274 225922 583342 225978
rect 583398 225922 583494 225978
rect 582874 208350 583494 225922
rect 582874 208294 582970 208350
rect 583026 208294 583094 208350
rect 583150 208294 583218 208350
rect 583274 208294 583342 208350
rect 583398 208294 583494 208350
rect 582874 208226 583494 208294
rect 582874 208170 582970 208226
rect 583026 208170 583094 208226
rect 583150 208170 583218 208226
rect 583274 208170 583342 208226
rect 583398 208170 583494 208226
rect 582874 208102 583494 208170
rect 582874 208046 582970 208102
rect 583026 208046 583094 208102
rect 583150 208046 583218 208102
rect 583274 208046 583342 208102
rect 583398 208046 583494 208102
rect 582874 207978 583494 208046
rect 582874 207922 582970 207978
rect 583026 207922 583094 207978
rect 583150 207922 583218 207978
rect 583274 207922 583342 207978
rect 583398 207922 583494 207978
rect 582874 190350 583494 207922
rect 582874 190294 582970 190350
rect 583026 190294 583094 190350
rect 583150 190294 583218 190350
rect 583274 190294 583342 190350
rect 583398 190294 583494 190350
rect 582874 190226 583494 190294
rect 582874 190170 582970 190226
rect 583026 190170 583094 190226
rect 583150 190170 583218 190226
rect 583274 190170 583342 190226
rect 583398 190170 583494 190226
rect 582874 190102 583494 190170
rect 582874 190046 582970 190102
rect 583026 190046 583094 190102
rect 583150 190046 583218 190102
rect 583274 190046 583342 190102
rect 583398 190046 583494 190102
rect 582874 189978 583494 190046
rect 582874 189922 582970 189978
rect 583026 189922 583094 189978
rect 583150 189922 583218 189978
rect 583274 189922 583342 189978
rect 583398 189922 583494 189978
rect 582874 172350 583494 189922
rect 582874 172294 582970 172350
rect 583026 172294 583094 172350
rect 583150 172294 583218 172350
rect 583274 172294 583342 172350
rect 583398 172294 583494 172350
rect 582874 172226 583494 172294
rect 582874 172170 582970 172226
rect 583026 172170 583094 172226
rect 583150 172170 583218 172226
rect 583274 172170 583342 172226
rect 583398 172170 583494 172226
rect 582874 172102 583494 172170
rect 582874 172046 582970 172102
rect 583026 172046 583094 172102
rect 583150 172046 583218 172102
rect 583274 172046 583342 172102
rect 583398 172046 583494 172102
rect 582874 171978 583494 172046
rect 582874 171922 582970 171978
rect 583026 171922 583094 171978
rect 583150 171922 583218 171978
rect 583274 171922 583342 171978
rect 583398 171922 583494 171978
rect 582874 154350 583494 171922
rect 582874 154294 582970 154350
rect 583026 154294 583094 154350
rect 583150 154294 583218 154350
rect 583274 154294 583342 154350
rect 583398 154294 583494 154350
rect 582874 154226 583494 154294
rect 582874 154170 582970 154226
rect 583026 154170 583094 154226
rect 583150 154170 583218 154226
rect 583274 154170 583342 154226
rect 583398 154170 583494 154226
rect 582874 154102 583494 154170
rect 582874 154046 582970 154102
rect 583026 154046 583094 154102
rect 583150 154046 583218 154102
rect 583274 154046 583342 154102
rect 583398 154046 583494 154102
rect 582874 153978 583494 154046
rect 582874 153922 582970 153978
rect 583026 153922 583094 153978
rect 583150 153922 583218 153978
rect 583274 153922 583342 153978
rect 583398 153922 583494 153978
rect 582874 136350 583494 153922
rect 582874 136294 582970 136350
rect 583026 136294 583094 136350
rect 583150 136294 583218 136350
rect 583274 136294 583342 136350
rect 583398 136294 583494 136350
rect 582874 136226 583494 136294
rect 582874 136170 582970 136226
rect 583026 136170 583094 136226
rect 583150 136170 583218 136226
rect 583274 136170 583342 136226
rect 583398 136170 583494 136226
rect 582874 136102 583494 136170
rect 582874 136046 582970 136102
rect 583026 136046 583094 136102
rect 583150 136046 583218 136102
rect 583274 136046 583342 136102
rect 583398 136046 583494 136102
rect 582874 135978 583494 136046
rect 582874 135922 582970 135978
rect 583026 135922 583094 135978
rect 583150 135922 583218 135978
rect 583274 135922 583342 135978
rect 583398 135922 583494 135978
rect 582874 118350 583494 135922
rect 582874 118294 582970 118350
rect 583026 118294 583094 118350
rect 583150 118294 583218 118350
rect 583274 118294 583342 118350
rect 583398 118294 583494 118350
rect 582874 118226 583494 118294
rect 582874 118170 582970 118226
rect 583026 118170 583094 118226
rect 583150 118170 583218 118226
rect 583274 118170 583342 118226
rect 583398 118170 583494 118226
rect 582874 118102 583494 118170
rect 582874 118046 582970 118102
rect 583026 118046 583094 118102
rect 583150 118046 583218 118102
rect 583274 118046 583342 118102
rect 583398 118046 583494 118102
rect 582874 117978 583494 118046
rect 582874 117922 582970 117978
rect 583026 117922 583094 117978
rect 583150 117922 583218 117978
rect 583274 117922 583342 117978
rect 583398 117922 583494 117978
rect 582874 100350 583494 117922
rect 582874 100294 582970 100350
rect 583026 100294 583094 100350
rect 583150 100294 583218 100350
rect 583274 100294 583342 100350
rect 583398 100294 583494 100350
rect 582874 100226 583494 100294
rect 582874 100170 582970 100226
rect 583026 100170 583094 100226
rect 583150 100170 583218 100226
rect 583274 100170 583342 100226
rect 583398 100170 583494 100226
rect 582874 100102 583494 100170
rect 582874 100046 582970 100102
rect 583026 100046 583094 100102
rect 583150 100046 583218 100102
rect 583274 100046 583342 100102
rect 583398 100046 583494 100102
rect 582874 99978 583494 100046
rect 582874 99922 582970 99978
rect 583026 99922 583094 99978
rect 583150 99922 583218 99978
rect 583274 99922 583342 99978
rect 583398 99922 583494 99978
rect 582874 82350 583494 99922
rect 582874 82294 582970 82350
rect 583026 82294 583094 82350
rect 583150 82294 583218 82350
rect 583274 82294 583342 82350
rect 583398 82294 583494 82350
rect 582874 82226 583494 82294
rect 582874 82170 582970 82226
rect 583026 82170 583094 82226
rect 583150 82170 583218 82226
rect 583274 82170 583342 82226
rect 583398 82170 583494 82226
rect 582874 82102 583494 82170
rect 582874 82046 582970 82102
rect 583026 82046 583094 82102
rect 583150 82046 583218 82102
rect 583274 82046 583342 82102
rect 583398 82046 583494 82102
rect 582874 81978 583494 82046
rect 582874 81922 582970 81978
rect 583026 81922 583094 81978
rect 583150 81922 583218 81978
rect 583274 81922 583342 81978
rect 583398 81922 583494 81978
rect 582874 64350 583494 81922
rect 582874 64294 582970 64350
rect 583026 64294 583094 64350
rect 583150 64294 583218 64350
rect 583274 64294 583342 64350
rect 583398 64294 583494 64350
rect 582874 64226 583494 64294
rect 582874 64170 582970 64226
rect 583026 64170 583094 64226
rect 583150 64170 583218 64226
rect 583274 64170 583342 64226
rect 583398 64170 583494 64226
rect 582874 64102 583494 64170
rect 582874 64046 582970 64102
rect 583026 64046 583094 64102
rect 583150 64046 583218 64102
rect 583274 64046 583342 64102
rect 583398 64046 583494 64102
rect 582874 63978 583494 64046
rect 582874 63922 582970 63978
rect 583026 63922 583094 63978
rect 583150 63922 583218 63978
rect 583274 63922 583342 63978
rect 583398 63922 583494 63978
rect 582874 46350 583494 63922
rect 582874 46294 582970 46350
rect 583026 46294 583094 46350
rect 583150 46294 583218 46350
rect 583274 46294 583342 46350
rect 583398 46294 583494 46350
rect 582874 46226 583494 46294
rect 582874 46170 582970 46226
rect 583026 46170 583094 46226
rect 583150 46170 583218 46226
rect 583274 46170 583342 46226
rect 583398 46170 583494 46226
rect 582874 46102 583494 46170
rect 582874 46046 582970 46102
rect 583026 46046 583094 46102
rect 583150 46046 583218 46102
rect 583274 46046 583342 46102
rect 583398 46046 583494 46102
rect 582874 45978 583494 46046
rect 582874 45922 582970 45978
rect 583026 45922 583094 45978
rect 583150 45922 583218 45978
rect 583274 45922 583342 45978
rect 583398 45922 583494 45978
rect 582874 28350 583494 45922
rect 582874 28294 582970 28350
rect 583026 28294 583094 28350
rect 583150 28294 583218 28350
rect 583274 28294 583342 28350
rect 583398 28294 583494 28350
rect 582874 28226 583494 28294
rect 582874 28170 582970 28226
rect 583026 28170 583094 28226
rect 583150 28170 583218 28226
rect 583274 28170 583342 28226
rect 583398 28170 583494 28226
rect 582874 28102 583494 28170
rect 582874 28046 582970 28102
rect 583026 28046 583094 28102
rect 583150 28046 583218 28102
rect 583274 28046 583342 28102
rect 583398 28046 583494 28102
rect 582874 27978 583494 28046
rect 582874 27922 582970 27978
rect 583026 27922 583094 27978
rect 583150 27922 583218 27978
rect 583274 27922 583342 27978
rect 583398 27922 583494 27978
rect 582874 10350 583494 27922
rect 582874 10294 582970 10350
rect 583026 10294 583094 10350
rect 583150 10294 583218 10350
rect 583274 10294 583342 10350
rect 583398 10294 583494 10350
rect 582874 10226 583494 10294
rect 582874 10170 582970 10226
rect 583026 10170 583094 10226
rect 583150 10170 583218 10226
rect 583274 10170 583342 10226
rect 583398 10170 583494 10226
rect 582874 10102 583494 10170
rect 582874 10046 582970 10102
rect 583026 10046 583094 10102
rect 583150 10046 583218 10102
rect 583274 10046 583342 10102
rect 583398 10046 583494 10102
rect 582874 9978 583494 10046
rect 582874 9922 582970 9978
rect 583026 9922 583094 9978
rect 583150 9922 583218 9978
rect 583274 9922 583342 9978
rect 583398 9922 583494 9978
rect 582874 -1120 583494 9922
rect 596400 597212 597020 597308
rect 596400 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect 596400 597088 597020 597156
rect 596400 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect 596400 596964 597020 597032
rect 596400 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect 596400 596840 597020 596908
rect 596400 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect 596400 580350 597020 596784
rect 596400 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597020 580350
rect 596400 580226 597020 580294
rect 596400 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597020 580226
rect 596400 580102 597020 580170
rect 596400 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597020 580102
rect 596400 579978 597020 580046
rect 596400 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597020 579978
rect 596400 562350 597020 579922
rect 596400 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597020 562350
rect 596400 562226 597020 562294
rect 596400 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597020 562226
rect 596400 562102 597020 562170
rect 596400 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597020 562102
rect 596400 561978 597020 562046
rect 596400 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597020 561978
rect 596400 544350 597020 561922
rect 596400 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597020 544350
rect 596400 544226 597020 544294
rect 596400 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597020 544226
rect 596400 544102 597020 544170
rect 596400 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597020 544102
rect 596400 543978 597020 544046
rect 596400 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597020 543978
rect 596400 526350 597020 543922
rect 596400 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597020 526350
rect 596400 526226 597020 526294
rect 596400 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597020 526226
rect 596400 526102 597020 526170
rect 596400 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597020 526102
rect 596400 525978 597020 526046
rect 596400 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597020 525978
rect 596400 508350 597020 525922
rect 596400 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597020 508350
rect 596400 508226 597020 508294
rect 596400 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597020 508226
rect 596400 508102 597020 508170
rect 596400 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597020 508102
rect 596400 507978 597020 508046
rect 596400 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597020 507978
rect 596400 490350 597020 507922
rect 596400 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597020 490350
rect 596400 490226 597020 490294
rect 596400 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597020 490226
rect 596400 490102 597020 490170
rect 596400 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597020 490102
rect 596400 489978 597020 490046
rect 596400 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597020 489978
rect 596400 472350 597020 489922
rect 596400 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597020 472350
rect 596400 472226 597020 472294
rect 596400 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597020 472226
rect 596400 472102 597020 472170
rect 596400 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597020 472102
rect 596400 471978 597020 472046
rect 596400 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597020 471978
rect 596400 454350 597020 471922
rect 596400 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597020 454350
rect 596400 454226 597020 454294
rect 596400 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597020 454226
rect 596400 454102 597020 454170
rect 596400 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597020 454102
rect 596400 453978 597020 454046
rect 596400 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597020 453978
rect 596400 436350 597020 453922
rect 596400 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597020 436350
rect 596400 436226 597020 436294
rect 596400 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597020 436226
rect 596400 436102 597020 436170
rect 596400 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597020 436102
rect 596400 435978 597020 436046
rect 596400 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597020 435978
rect 596400 418350 597020 435922
rect 596400 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597020 418350
rect 596400 418226 597020 418294
rect 596400 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597020 418226
rect 596400 418102 597020 418170
rect 596400 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597020 418102
rect 596400 417978 597020 418046
rect 596400 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597020 417978
rect 596400 400350 597020 417922
rect 596400 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597020 400350
rect 596400 400226 597020 400294
rect 596400 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597020 400226
rect 596400 400102 597020 400170
rect 596400 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597020 400102
rect 596400 399978 597020 400046
rect 596400 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597020 399978
rect 596400 382350 597020 399922
rect 596400 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597020 382350
rect 596400 382226 597020 382294
rect 596400 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597020 382226
rect 596400 382102 597020 382170
rect 596400 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597020 382102
rect 596400 381978 597020 382046
rect 596400 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597020 381978
rect 596400 364350 597020 381922
rect 596400 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597020 364350
rect 596400 364226 597020 364294
rect 596400 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597020 364226
rect 596400 364102 597020 364170
rect 596400 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597020 364102
rect 596400 363978 597020 364046
rect 596400 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597020 363978
rect 596400 346350 597020 363922
rect 596400 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597020 346350
rect 596400 346226 597020 346294
rect 596400 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597020 346226
rect 596400 346102 597020 346170
rect 596400 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597020 346102
rect 596400 345978 597020 346046
rect 596400 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597020 345978
rect 596400 328350 597020 345922
rect 596400 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597020 328350
rect 596400 328226 597020 328294
rect 596400 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597020 328226
rect 596400 328102 597020 328170
rect 596400 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597020 328102
rect 596400 327978 597020 328046
rect 596400 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597020 327978
rect 596400 310350 597020 327922
rect 596400 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597020 310350
rect 596400 310226 597020 310294
rect 596400 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597020 310226
rect 596400 310102 597020 310170
rect 596400 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597020 310102
rect 596400 309978 597020 310046
rect 596400 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597020 309978
rect 596400 292350 597020 309922
rect 596400 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597020 292350
rect 596400 292226 597020 292294
rect 596400 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597020 292226
rect 596400 292102 597020 292170
rect 596400 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597020 292102
rect 596400 291978 597020 292046
rect 596400 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597020 291978
rect 596400 274350 597020 291922
rect 596400 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597020 274350
rect 596400 274226 597020 274294
rect 596400 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597020 274226
rect 596400 274102 597020 274170
rect 596400 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597020 274102
rect 596400 273978 597020 274046
rect 596400 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597020 273978
rect 596400 256350 597020 273922
rect 596400 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597020 256350
rect 596400 256226 597020 256294
rect 596400 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597020 256226
rect 596400 256102 597020 256170
rect 596400 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597020 256102
rect 596400 255978 597020 256046
rect 596400 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597020 255978
rect 596400 238350 597020 255922
rect 596400 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597020 238350
rect 596400 238226 597020 238294
rect 596400 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597020 238226
rect 596400 238102 597020 238170
rect 596400 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597020 238102
rect 596400 237978 597020 238046
rect 596400 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597020 237978
rect 596400 220350 597020 237922
rect 596400 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597020 220350
rect 596400 220226 597020 220294
rect 596400 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597020 220226
rect 596400 220102 597020 220170
rect 596400 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597020 220102
rect 596400 219978 597020 220046
rect 596400 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597020 219978
rect 596400 202350 597020 219922
rect 596400 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597020 202350
rect 596400 202226 597020 202294
rect 596400 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597020 202226
rect 596400 202102 597020 202170
rect 596400 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597020 202102
rect 596400 201978 597020 202046
rect 596400 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597020 201978
rect 596400 184350 597020 201922
rect 596400 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597020 184350
rect 596400 184226 597020 184294
rect 596400 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597020 184226
rect 596400 184102 597020 184170
rect 596400 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597020 184102
rect 596400 183978 597020 184046
rect 596400 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597020 183978
rect 596400 166350 597020 183922
rect 596400 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597020 166350
rect 596400 166226 597020 166294
rect 596400 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597020 166226
rect 596400 166102 597020 166170
rect 596400 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597020 166102
rect 596400 165978 597020 166046
rect 596400 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597020 165978
rect 596400 148350 597020 165922
rect 596400 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597020 148350
rect 596400 148226 597020 148294
rect 596400 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597020 148226
rect 596400 148102 597020 148170
rect 596400 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597020 148102
rect 596400 147978 597020 148046
rect 596400 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597020 147978
rect 596400 130350 597020 147922
rect 596400 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597020 130350
rect 596400 130226 597020 130294
rect 596400 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597020 130226
rect 596400 130102 597020 130170
rect 596400 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597020 130102
rect 596400 129978 597020 130046
rect 596400 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597020 129978
rect 596400 112350 597020 129922
rect 596400 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597020 112350
rect 596400 112226 597020 112294
rect 596400 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597020 112226
rect 596400 112102 597020 112170
rect 596400 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597020 112102
rect 596400 111978 597020 112046
rect 596400 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597020 111978
rect 596400 94350 597020 111922
rect 596400 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597020 94350
rect 596400 94226 597020 94294
rect 596400 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597020 94226
rect 596400 94102 597020 94170
rect 596400 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597020 94102
rect 596400 93978 597020 94046
rect 596400 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597020 93978
rect 596400 76350 597020 93922
rect 596400 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597020 76350
rect 596400 76226 597020 76294
rect 596400 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597020 76226
rect 596400 76102 597020 76170
rect 596400 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597020 76102
rect 596400 75978 597020 76046
rect 596400 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597020 75978
rect 596400 58350 597020 75922
rect 596400 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597020 58350
rect 596400 58226 597020 58294
rect 596400 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597020 58226
rect 596400 58102 597020 58170
rect 596400 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597020 58102
rect 596400 57978 597020 58046
rect 596400 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597020 57978
rect 596400 40350 597020 57922
rect 596400 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597020 40350
rect 596400 40226 597020 40294
rect 596400 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597020 40226
rect 596400 40102 597020 40170
rect 596400 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597020 40102
rect 596400 39978 597020 40046
rect 596400 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597020 39978
rect 596400 22350 597020 39922
rect 596400 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597020 22350
rect 596400 22226 597020 22294
rect 596400 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597020 22226
rect 596400 22102 597020 22170
rect 596400 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597020 22102
rect 596400 21978 597020 22046
rect 596400 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597020 21978
rect 596400 4350 597020 21922
rect 596400 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597020 4350
rect 596400 4226 597020 4294
rect 596400 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597020 4226
rect 596400 4102 597020 4170
rect 596400 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597020 4102
rect 596400 3978 597020 4046
rect 596400 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597020 3978
rect 596400 -160 597020 3922
rect 596400 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect 596400 -284 597020 -216
rect 596400 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect 596400 -408 597020 -340
rect 596400 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect 596400 -532 597020 -464
rect 596400 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect 596400 -684 597020 -588
rect 597360 586350 597980 597744
rect 597360 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect 597360 586226 597980 586294
rect 597360 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect 597360 586102 597980 586170
rect 597360 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect 597360 585978 597980 586046
rect 597360 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect 597360 568350 597980 585922
rect 597360 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect 597360 568226 597980 568294
rect 597360 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect 597360 568102 597980 568170
rect 597360 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect 597360 567978 597980 568046
rect 597360 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect 597360 550350 597980 567922
rect 597360 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect 597360 550226 597980 550294
rect 597360 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect 597360 550102 597980 550170
rect 597360 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect 597360 549978 597980 550046
rect 597360 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect 597360 532350 597980 549922
rect 597360 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect 597360 532226 597980 532294
rect 597360 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect 597360 532102 597980 532170
rect 597360 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect 597360 531978 597980 532046
rect 597360 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect 597360 514350 597980 531922
rect 597360 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect 597360 514226 597980 514294
rect 597360 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect 597360 514102 597980 514170
rect 597360 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect 597360 513978 597980 514046
rect 597360 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect 597360 496350 597980 513922
rect 597360 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect 597360 496226 597980 496294
rect 597360 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect 597360 496102 597980 496170
rect 597360 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect 597360 495978 597980 496046
rect 597360 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect 597360 478350 597980 495922
rect 597360 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect 597360 478226 597980 478294
rect 597360 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect 597360 478102 597980 478170
rect 597360 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect 597360 477978 597980 478046
rect 597360 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect 597360 460350 597980 477922
rect 597360 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect 597360 460226 597980 460294
rect 597360 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect 597360 460102 597980 460170
rect 597360 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect 597360 459978 597980 460046
rect 597360 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect 597360 442350 597980 459922
rect 597360 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect 597360 442226 597980 442294
rect 597360 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect 597360 442102 597980 442170
rect 597360 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect 597360 441978 597980 442046
rect 597360 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect 597360 424350 597980 441922
rect 597360 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect 597360 424226 597980 424294
rect 597360 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect 597360 424102 597980 424170
rect 597360 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect 597360 423978 597980 424046
rect 597360 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect 597360 406350 597980 423922
rect 597360 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect 597360 406226 597980 406294
rect 597360 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect 597360 406102 597980 406170
rect 597360 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect 597360 405978 597980 406046
rect 597360 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect 597360 388350 597980 405922
rect 597360 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect 597360 388226 597980 388294
rect 597360 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect 597360 388102 597980 388170
rect 597360 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect 597360 387978 597980 388046
rect 597360 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect 597360 370350 597980 387922
rect 597360 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect 597360 370226 597980 370294
rect 597360 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect 597360 370102 597980 370170
rect 597360 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect 597360 369978 597980 370046
rect 597360 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect 597360 352350 597980 369922
rect 597360 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect 597360 352226 597980 352294
rect 597360 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect 597360 352102 597980 352170
rect 597360 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect 597360 351978 597980 352046
rect 597360 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect 597360 334350 597980 351922
rect 597360 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect 597360 334226 597980 334294
rect 597360 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect 597360 334102 597980 334170
rect 597360 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect 597360 333978 597980 334046
rect 597360 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect 597360 316350 597980 333922
rect 597360 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect 597360 316226 597980 316294
rect 597360 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect 597360 316102 597980 316170
rect 597360 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect 597360 315978 597980 316046
rect 597360 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect 597360 298350 597980 315922
rect 597360 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect 597360 298226 597980 298294
rect 597360 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect 597360 298102 597980 298170
rect 597360 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect 597360 297978 597980 298046
rect 597360 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect 597360 280350 597980 297922
rect 597360 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect 597360 280226 597980 280294
rect 597360 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect 597360 280102 597980 280170
rect 597360 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect 597360 279978 597980 280046
rect 597360 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect 597360 262350 597980 279922
rect 597360 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect 597360 262226 597980 262294
rect 597360 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect 597360 262102 597980 262170
rect 597360 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect 597360 261978 597980 262046
rect 597360 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect 597360 244350 597980 261922
rect 597360 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect 597360 244226 597980 244294
rect 597360 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect 597360 244102 597980 244170
rect 597360 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect 597360 243978 597980 244046
rect 597360 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect 597360 226350 597980 243922
rect 597360 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect 597360 226226 597980 226294
rect 597360 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect 597360 226102 597980 226170
rect 597360 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect 597360 225978 597980 226046
rect 597360 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect 597360 208350 597980 225922
rect 597360 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect 597360 208226 597980 208294
rect 597360 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect 597360 208102 597980 208170
rect 597360 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect 597360 207978 597980 208046
rect 597360 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect 597360 190350 597980 207922
rect 597360 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect 597360 190226 597980 190294
rect 597360 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect 597360 190102 597980 190170
rect 597360 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect 597360 189978 597980 190046
rect 597360 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect 597360 172350 597980 189922
rect 597360 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect 597360 172226 597980 172294
rect 597360 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect 597360 172102 597980 172170
rect 597360 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect 597360 171978 597980 172046
rect 597360 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect 597360 154350 597980 171922
rect 597360 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect 597360 154226 597980 154294
rect 597360 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect 597360 154102 597980 154170
rect 597360 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect 597360 153978 597980 154046
rect 597360 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect 597360 136350 597980 153922
rect 597360 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect 597360 136226 597980 136294
rect 597360 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect 597360 136102 597980 136170
rect 597360 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect 597360 135978 597980 136046
rect 597360 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect 597360 118350 597980 135922
rect 597360 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect 597360 118226 597980 118294
rect 597360 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect 597360 118102 597980 118170
rect 597360 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect 597360 117978 597980 118046
rect 597360 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect 597360 100350 597980 117922
rect 597360 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect 597360 100226 597980 100294
rect 597360 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect 597360 100102 597980 100170
rect 597360 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect 597360 99978 597980 100046
rect 597360 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect 597360 82350 597980 99922
rect 597360 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect 597360 82226 597980 82294
rect 597360 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect 597360 82102 597980 82170
rect 597360 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect 597360 81978 597980 82046
rect 597360 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect 597360 64350 597980 81922
rect 597360 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect 597360 64226 597980 64294
rect 597360 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect 597360 64102 597980 64170
rect 597360 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect 597360 63978 597980 64046
rect 597360 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect 597360 46350 597980 63922
rect 597360 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect 597360 46226 597980 46294
rect 597360 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect 597360 46102 597980 46170
rect 597360 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect 597360 45978 597980 46046
rect 597360 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect 597360 28350 597980 45922
rect 597360 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect 597360 28226 597980 28294
rect 597360 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect 597360 28102 597980 28170
rect 597360 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect 597360 27978 597980 28046
rect 597360 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect 597360 10350 597980 27922
rect 597360 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect 597360 10226 597980 10294
rect 597360 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect 597360 10102 597980 10170
rect 597360 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect 597360 9978 597980 10046
rect 597360 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect 582874 -1176 582970 -1120
rect 583026 -1176 583094 -1120
rect 583150 -1176 583218 -1120
rect 583274 -1176 583342 -1120
rect 583398 -1176 583494 -1120
rect 582874 -1244 583494 -1176
rect 582874 -1300 582970 -1244
rect 583026 -1300 583094 -1244
rect 583150 -1300 583218 -1244
rect 583274 -1300 583342 -1244
rect 583398 -1300 583494 -1244
rect 582874 -1368 583494 -1300
rect 582874 -1424 582970 -1368
rect 583026 -1424 583094 -1368
rect 583150 -1424 583218 -1368
rect 583274 -1424 583342 -1368
rect 583398 -1424 583494 -1368
rect 582874 -1492 583494 -1424
rect 582874 -1548 582970 -1492
rect 583026 -1548 583094 -1492
rect 583150 -1548 583218 -1492
rect 583274 -1548 583342 -1492
rect 583398 -1548 583494 -1492
rect 582874 -1644 583494 -1548
rect 597360 -1120 597980 9922
rect 597360 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect 597360 -1244 597980 -1176
rect 597360 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect 597360 -1368 597980 -1300
rect 597360 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect 597360 -1492 597980 -1424
rect 597360 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect 597360 -1644 597980 -1548
<< via4 >>
rect -1820 598116 -1764 598172
rect -1696 598116 -1640 598172
rect -1572 598116 -1516 598172
rect -1448 598116 -1392 598172
rect -1820 597992 -1764 598048
rect -1696 597992 -1640 598048
rect -1572 597992 -1516 598048
rect -1448 597992 -1392 598048
rect -1820 597868 -1764 597924
rect -1696 597868 -1640 597924
rect -1572 597868 -1516 597924
rect -1448 597868 -1392 597924
rect -1820 597744 -1764 597800
rect -1696 597744 -1640 597800
rect -1572 597744 -1516 597800
rect -1448 597744 -1392 597800
rect -1820 586294 -1764 586350
rect -1696 586294 -1640 586350
rect -1572 586294 -1516 586350
rect -1448 586294 -1392 586350
rect -1820 586170 -1764 586226
rect -1696 586170 -1640 586226
rect -1572 586170 -1516 586226
rect -1448 586170 -1392 586226
rect -1820 586046 -1764 586102
rect -1696 586046 -1640 586102
rect -1572 586046 -1516 586102
rect -1448 586046 -1392 586102
rect -1820 585922 -1764 585978
rect -1696 585922 -1640 585978
rect -1572 585922 -1516 585978
rect -1448 585922 -1392 585978
rect -1820 568294 -1764 568350
rect -1696 568294 -1640 568350
rect -1572 568294 -1516 568350
rect -1448 568294 -1392 568350
rect -1820 568170 -1764 568226
rect -1696 568170 -1640 568226
rect -1572 568170 -1516 568226
rect -1448 568170 -1392 568226
rect -1820 568046 -1764 568102
rect -1696 568046 -1640 568102
rect -1572 568046 -1516 568102
rect -1448 568046 -1392 568102
rect -1820 567922 -1764 567978
rect -1696 567922 -1640 567978
rect -1572 567922 -1516 567978
rect -1448 567922 -1392 567978
rect -1820 550294 -1764 550350
rect -1696 550294 -1640 550350
rect -1572 550294 -1516 550350
rect -1448 550294 -1392 550350
rect -1820 550170 -1764 550226
rect -1696 550170 -1640 550226
rect -1572 550170 -1516 550226
rect -1448 550170 -1392 550226
rect -1820 550046 -1764 550102
rect -1696 550046 -1640 550102
rect -1572 550046 -1516 550102
rect -1448 550046 -1392 550102
rect -1820 549922 -1764 549978
rect -1696 549922 -1640 549978
rect -1572 549922 -1516 549978
rect -1448 549922 -1392 549978
rect -1820 532294 -1764 532350
rect -1696 532294 -1640 532350
rect -1572 532294 -1516 532350
rect -1448 532294 -1392 532350
rect -1820 532170 -1764 532226
rect -1696 532170 -1640 532226
rect -1572 532170 -1516 532226
rect -1448 532170 -1392 532226
rect -1820 532046 -1764 532102
rect -1696 532046 -1640 532102
rect -1572 532046 -1516 532102
rect -1448 532046 -1392 532102
rect -1820 531922 -1764 531978
rect -1696 531922 -1640 531978
rect -1572 531922 -1516 531978
rect -1448 531922 -1392 531978
rect -1820 514294 -1764 514350
rect -1696 514294 -1640 514350
rect -1572 514294 -1516 514350
rect -1448 514294 -1392 514350
rect -1820 514170 -1764 514226
rect -1696 514170 -1640 514226
rect -1572 514170 -1516 514226
rect -1448 514170 -1392 514226
rect -1820 514046 -1764 514102
rect -1696 514046 -1640 514102
rect -1572 514046 -1516 514102
rect -1448 514046 -1392 514102
rect -1820 513922 -1764 513978
rect -1696 513922 -1640 513978
rect -1572 513922 -1516 513978
rect -1448 513922 -1392 513978
rect -1820 496294 -1764 496350
rect -1696 496294 -1640 496350
rect -1572 496294 -1516 496350
rect -1448 496294 -1392 496350
rect -1820 496170 -1764 496226
rect -1696 496170 -1640 496226
rect -1572 496170 -1516 496226
rect -1448 496170 -1392 496226
rect -1820 496046 -1764 496102
rect -1696 496046 -1640 496102
rect -1572 496046 -1516 496102
rect -1448 496046 -1392 496102
rect -1820 495922 -1764 495978
rect -1696 495922 -1640 495978
rect -1572 495922 -1516 495978
rect -1448 495922 -1392 495978
rect -1820 478294 -1764 478350
rect -1696 478294 -1640 478350
rect -1572 478294 -1516 478350
rect -1448 478294 -1392 478350
rect -1820 478170 -1764 478226
rect -1696 478170 -1640 478226
rect -1572 478170 -1516 478226
rect -1448 478170 -1392 478226
rect -1820 478046 -1764 478102
rect -1696 478046 -1640 478102
rect -1572 478046 -1516 478102
rect -1448 478046 -1392 478102
rect -1820 477922 -1764 477978
rect -1696 477922 -1640 477978
rect -1572 477922 -1516 477978
rect -1448 477922 -1392 477978
rect -1820 460294 -1764 460350
rect -1696 460294 -1640 460350
rect -1572 460294 -1516 460350
rect -1448 460294 -1392 460350
rect -1820 460170 -1764 460226
rect -1696 460170 -1640 460226
rect -1572 460170 -1516 460226
rect -1448 460170 -1392 460226
rect -1820 460046 -1764 460102
rect -1696 460046 -1640 460102
rect -1572 460046 -1516 460102
rect -1448 460046 -1392 460102
rect -1820 459922 -1764 459978
rect -1696 459922 -1640 459978
rect -1572 459922 -1516 459978
rect -1448 459922 -1392 459978
rect -1820 442294 -1764 442350
rect -1696 442294 -1640 442350
rect -1572 442294 -1516 442350
rect -1448 442294 -1392 442350
rect -1820 442170 -1764 442226
rect -1696 442170 -1640 442226
rect -1572 442170 -1516 442226
rect -1448 442170 -1392 442226
rect -1820 442046 -1764 442102
rect -1696 442046 -1640 442102
rect -1572 442046 -1516 442102
rect -1448 442046 -1392 442102
rect -1820 441922 -1764 441978
rect -1696 441922 -1640 441978
rect -1572 441922 -1516 441978
rect -1448 441922 -1392 441978
rect -1820 424294 -1764 424350
rect -1696 424294 -1640 424350
rect -1572 424294 -1516 424350
rect -1448 424294 -1392 424350
rect -1820 424170 -1764 424226
rect -1696 424170 -1640 424226
rect -1572 424170 -1516 424226
rect -1448 424170 -1392 424226
rect -1820 424046 -1764 424102
rect -1696 424046 -1640 424102
rect -1572 424046 -1516 424102
rect -1448 424046 -1392 424102
rect -1820 423922 -1764 423978
rect -1696 423922 -1640 423978
rect -1572 423922 -1516 423978
rect -1448 423922 -1392 423978
rect -1820 406294 -1764 406350
rect -1696 406294 -1640 406350
rect -1572 406294 -1516 406350
rect -1448 406294 -1392 406350
rect -1820 406170 -1764 406226
rect -1696 406170 -1640 406226
rect -1572 406170 -1516 406226
rect -1448 406170 -1392 406226
rect -1820 406046 -1764 406102
rect -1696 406046 -1640 406102
rect -1572 406046 -1516 406102
rect -1448 406046 -1392 406102
rect -1820 405922 -1764 405978
rect -1696 405922 -1640 405978
rect -1572 405922 -1516 405978
rect -1448 405922 -1392 405978
rect -1820 388294 -1764 388350
rect -1696 388294 -1640 388350
rect -1572 388294 -1516 388350
rect -1448 388294 -1392 388350
rect -1820 388170 -1764 388226
rect -1696 388170 -1640 388226
rect -1572 388170 -1516 388226
rect -1448 388170 -1392 388226
rect -1820 388046 -1764 388102
rect -1696 388046 -1640 388102
rect -1572 388046 -1516 388102
rect -1448 388046 -1392 388102
rect -1820 387922 -1764 387978
rect -1696 387922 -1640 387978
rect -1572 387922 -1516 387978
rect -1448 387922 -1392 387978
rect -1820 370294 -1764 370350
rect -1696 370294 -1640 370350
rect -1572 370294 -1516 370350
rect -1448 370294 -1392 370350
rect -1820 370170 -1764 370226
rect -1696 370170 -1640 370226
rect -1572 370170 -1516 370226
rect -1448 370170 -1392 370226
rect -1820 370046 -1764 370102
rect -1696 370046 -1640 370102
rect -1572 370046 -1516 370102
rect -1448 370046 -1392 370102
rect -1820 369922 -1764 369978
rect -1696 369922 -1640 369978
rect -1572 369922 -1516 369978
rect -1448 369922 -1392 369978
rect -1820 352294 -1764 352350
rect -1696 352294 -1640 352350
rect -1572 352294 -1516 352350
rect -1448 352294 -1392 352350
rect -1820 352170 -1764 352226
rect -1696 352170 -1640 352226
rect -1572 352170 -1516 352226
rect -1448 352170 -1392 352226
rect -1820 352046 -1764 352102
rect -1696 352046 -1640 352102
rect -1572 352046 -1516 352102
rect -1448 352046 -1392 352102
rect -1820 351922 -1764 351978
rect -1696 351922 -1640 351978
rect -1572 351922 -1516 351978
rect -1448 351922 -1392 351978
rect -1820 334294 -1764 334350
rect -1696 334294 -1640 334350
rect -1572 334294 -1516 334350
rect -1448 334294 -1392 334350
rect -1820 334170 -1764 334226
rect -1696 334170 -1640 334226
rect -1572 334170 -1516 334226
rect -1448 334170 -1392 334226
rect -1820 334046 -1764 334102
rect -1696 334046 -1640 334102
rect -1572 334046 -1516 334102
rect -1448 334046 -1392 334102
rect -1820 333922 -1764 333978
rect -1696 333922 -1640 333978
rect -1572 333922 -1516 333978
rect -1448 333922 -1392 333978
rect -1820 316294 -1764 316350
rect -1696 316294 -1640 316350
rect -1572 316294 -1516 316350
rect -1448 316294 -1392 316350
rect -1820 316170 -1764 316226
rect -1696 316170 -1640 316226
rect -1572 316170 -1516 316226
rect -1448 316170 -1392 316226
rect -1820 316046 -1764 316102
rect -1696 316046 -1640 316102
rect -1572 316046 -1516 316102
rect -1448 316046 -1392 316102
rect -1820 315922 -1764 315978
rect -1696 315922 -1640 315978
rect -1572 315922 -1516 315978
rect -1448 315922 -1392 315978
rect -1820 298294 -1764 298350
rect -1696 298294 -1640 298350
rect -1572 298294 -1516 298350
rect -1448 298294 -1392 298350
rect -1820 298170 -1764 298226
rect -1696 298170 -1640 298226
rect -1572 298170 -1516 298226
rect -1448 298170 -1392 298226
rect -1820 298046 -1764 298102
rect -1696 298046 -1640 298102
rect -1572 298046 -1516 298102
rect -1448 298046 -1392 298102
rect -1820 297922 -1764 297978
rect -1696 297922 -1640 297978
rect -1572 297922 -1516 297978
rect -1448 297922 -1392 297978
rect -1820 280294 -1764 280350
rect -1696 280294 -1640 280350
rect -1572 280294 -1516 280350
rect -1448 280294 -1392 280350
rect -1820 280170 -1764 280226
rect -1696 280170 -1640 280226
rect -1572 280170 -1516 280226
rect -1448 280170 -1392 280226
rect -1820 280046 -1764 280102
rect -1696 280046 -1640 280102
rect -1572 280046 -1516 280102
rect -1448 280046 -1392 280102
rect -1820 279922 -1764 279978
rect -1696 279922 -1640 279978
rect -1572 279922 -1516 279978
rect -1448 279922 -1392 279978
rect -1820 262294 -1764 262350
rect -1696 262294 -1640 262350
rect -1572 262294 -1516 262350
rect -1448 262294 -1392 262350
rect -1820 262170 -1764 262226
rect -1696 262170 -1640 262226
rect -1572 262170 -1516 262226
rect -1448 262170 -1392 262226
rect -1820 262046 -1764 262102
rect -1696 262046 -1640 262102
rect -1572 262046 -1516 262102
rect -1448 262046 -1392 262102
rect -1820 261922 -1764 261978
rect -1696 261922 -1640 261978
rect -1572 261922 -1516 261978
rect -1448 261922 -1392 261978
rect -1820 244294 -1764 244350
rect -1696 244294 -1640 244350
rect -1572 244294 -1516 244350
rect -1448 244294 -1392 244350
rect -1820 244170 -1764 244226
rect -1696 244170 -1640 244226
rect -1572 244170 -1516 244226
rect -1448 244170 -1392 244226
rect -1820 244046 -1764 244102
rect -1696 244046 -1640 244102
rect -1572 244046 -1516 244102
rect -1448 244046 -1392 244102
rect -1820 243922 -1764 243978
rect -1696 243922 -1640 243978
rect -1572 243922 -1516 243978
rect -1448 243922 -1392 243978
rect -1820 226294 -1764 226350
rect -1696 226294 -1640 226350
rect -1572 226294 -1516 226350
rect -1448 226294 -1392 226350
rect -1820 226170 -1764 226226
rect -1696 226170 -1640 226226
rect -1572 226170 -1516 226226
rect -1448 226170 -1392 226226
rect -1820 226046 -1764 226102
rect -1696 226046 -1640 226102
rect -1572 226046 -1516 226102
rect -1448 226046 -1392 226102
rect -1820 225922 -1764 225978
rect -1696 225922 -1640 225978
rect -1572 225922 -1516 225978
rect -1448 225922 -1392 225978
rect -1820 208294 -1764 208350
rect -1696 208294 -1640 208350
rect -1572 208294 -1516 208350
rect -1448 208294 -1392 208350
rect -1820 208170 -1764 208226
rect -1696 208170 -1640 208226
rect -1572 208170 -1516 208226
rect -1448 208170 -1392 208226
rect -1820 208046 -1764 208102
rect -1696 208046 -1640 208102
rect -1572 208046 -1516 208102
rect -1448 208046 -1392 208102
rect -1820 207922 -1764 207978
rect -1696 207922 -1640 207978
rect -1572 207922 -1516 207978
rect -1448 207922 -1392 207978
rect -1820 190294 -1764 190350
rect -1696 190294 -1640 190350
rect -1572 190294 -1516 190350
rect -1448 190294 -1392 190350
rect -1820 190170 -1764 190226
rect -1696 190170 -1640 190226
rect -1572 190170 -1516 190226
rect -1448 190170 -1392 190226
rect -1820 190046 -1764 190102
rect -1696 190046 -1640 190102
rect -1572 190046 -1516 190102
rect -1448 190046 -1392 190102
rect -1820 189922 -1764 189978
rect -1696 189922 -1640 189978
rect -1572 189922 -1516 189978
rect -1448 189922 -1392 189978
rect -1820 172294 -1764 172350
rect -1696 172294 -1640 172350
rect -1572 172294 -1516 172350
rect -1448 172294 -1392 172350
rect -1820 172170 -1764 172226
rect -1696 172170 -1640 172226
rect -1572 172170 -1516 172226
rect -1448 172170 -1392 172226
rect -1820 172046 -1764 172102
rect -1696 172046 -1640 172102
rect -1572 172046 -1516 172102
rect -1448 172046 -1392 172102
rect -1820 171922 -1764 171978
rect -1696 171922 -1640 171978
rect -1572 171922 -1516 171978
rect -1448 171922 -1392 171978
rect -1820 154294 -1764 154350
rect -1696 154294 -1640 154350
rect -1572 154294 -1516 154350
rect -1448 154294 -1392 154350
rect -1820 154170 -1764 154226
rect -1696 154170 -1640 154226
rect -1572 154170 -1516 154226
rect -1448 154170 -1392 154226
rect -1820 154046 -1764 154102
rect -1696 154046 -1640 154102
rect -1572 154046 -1516 154102
rect -1448 154046 -1392 154102
rect -1820 153922 -1764 153978
rect -1696 153922 -1640 153978
rect -1572 153922 -1516 153978
rect -1448 153922 -1392 153978
rect -1820 136294 -1764 136350
rect -1696 136294 -1640 136350
rect -1572 136294 -1516 136350
rect -1448 136294 -1392 136350
rect -1820 136170 -1764 136226
rect -1696 136170 -1640 136226
rect -1572 136170 -1516 136226
rect -1448 136170 -1392 136226
rect -1820 136046 -1764 136102
rect -1696 136046 -1640 136102
rect -1572 136046 -1516 136102
rect -1448 136046 -1392 136102
rect -1820 135922 -1764 135978
rect -1696 135922 -1640 135978
rect -1572 135922 -1516 135978
rect -1448 135922 -1392 135978
rect -1820 118294 -1764 118350
rect -1696 118294 -1640 118350
rect -1572 118294 -1516 118350
rect -1448 118294 -1392 118350
rect -1820 118170 -1764 118226
rect -1696 118170 -1640 118226
rect -1572 118170 -1516 118226
rect -1448 118170 -1392 118226
rect -1820 118046 -1764 118102
rect -1696 118046 -1640 118102
rect -1572 118046 -1516 118102
rect -1448 118046 -1392 118102
rect -1820 117922 -1764 117978
rect -1696 117922 -1640 117978
rect -1572 117922 -1516 117978
rect -1448 117922 -1392 117978
rect -1820 100294 -1764 100350
rect -1696 100294 -1640 100350
rect -1572 100294 -1516 100350
rect -1448 100294 -1392 100350
rect -1820 100170 -1764 100226
rect -1696 100170 -1640 100226
rect -1572 100170 -1516 100226
rect -1448 100170 -1392 100226
rect -1820 100046 -1764 100102
rect -1696 100046 -1640 100102
rect -1572 100046 -1516 100102
rect -1448 100046 -1392 100102
rect -1820 99922 -1764 99978
rect -1696 99922 -1640 99978
rect -1572 99922 -1516 99978
rect -1448 99922 -1392 99978
rect -1820 82294 -1764 82350
rect -1696 82294 -1640 82350
rect -1572 82294 -1516 82350
rect -1448 82294 -1392 82350
rect -1820 82170 -1764 82226
rect -1696 82170 -1640 82226
rect -1572 82170 -1516 82226
rect -1448 82170 -1392 82226
rect -1820 82046 -1764 82102
rect -1696 82046 -1640 82102
rect -1572 82046 -1516 82102
rect -1448 82046 -1392 82102
rect -1820 81922 -1764 81978
rect -1696 81922 -1640 81978
rect -1572 81922 -1516 81978
rect -1448 81922 -1392 81978
rect -1820 64294 -1764 64350
rect -1696 64294 -1640 64350
rect -1572 64294 -1516 64350
rect -1448 64294 -1392 64350
rect -1820 64170 -1764 64226
rect -1696 64170 -1640 64226
rect -1572 64170 -1516 64226
rect -1448 64170 -1392 64226
rect -1820 64046 -1764 64102
rect -1696 64046 -1640 64102
rect -1572 64046 -1516 64102
rect -1448 64046 -1392 64102
rect -1820 63922 -1764 63978
rect -1696 63922 -1640 63978
rect -1572 63922 -1516 63978
rect -1448 63922 -1392 63978
rect -1820 46294 -1764 46350
rect -1696 46294 -1640 46350
rect -1572 46294 -1516 46350
rect -1448 46294 -1392 46350
rect -1820 46170 -1764 46226
rect -1696 46170 -1640 46226
rect -1572 46170 -1516 46226
rect -1448 46170 -1392 46226
rect -1820 46046 -1764 46102
rect -1696 46046 -1640 46102
rect -1572 46046 -1516 46102
rect -1448 46046 -1392 46102
rect -1820 45922 -1764 45978
rect -1696 45922 -1640 45978
rect -1572 45922 -1516 45978
rect -1448 45922 -1392 45978
rect -1820 28294 -1764 28350
rect -1696 28294 -1640 28350
rect -1572 28294 -1516 28350
rect -1448 28294 -1392 28350
rect -1820 28170 -1764 28226
rect -1696 28170 -1640 28226
rect -1572 28170 -1516 28226
rect -1448 28170 -1392 28226
rect -1820 28046 -1764 28102
rect -1696 28046 -1640 28102
rect -1572 28046 -1516 28102
rect -1448 28046 -1392 28102
rect -1820 27922 -1764 27978
rect -1696 27922 -1640 27978
rect -1572 27922 -1516 27978
rect -1448 27922 -1392 27978
rect -1820 10294 -1764 10350
rect -1696 10294 -1640 10350
rect -1572 10294 -1516 10350
rect -1448 10294 -1392 10350
rect -1820 10170 -1764 10226
rect -1696 10170 -1640 10226
rect -1572 10170 -1516 10226
rect -1448 10170 -1392 10226
rect -1820 10046 -1764 10102
rect -1696 10046 -1640 10102
rect -1572 10046 -1516 10102
rect -1448 10046 -1392 10102
rect -1820 9922 -1764 9978
rect -1696 9922 -1640 9978
rect -1572 9922 -1516 9978
rect -1448 9922 -1392 9978
rect -860 597156 -804 597212
rect -736 597156 -680 597212
rect -612 597156 -556 597212
rect -488 597156 -432 597212
rect -860 597032 -804 597088
rect -736 597032 -680 597088
rect -612 597032 -556 597088
rect -488 597032 -432 597088
rect -860 596908 -804 596964
rect -736 596908 -680 596964
rect -612 596908 -556 596964
rect -488 596908 -432 596964
rect -860 596784 -804 596840
rect -736 596784 -680 596840
rect -612 596784 -556 596840
rect -488 596784 -432 596840
rect -860 580294 -804 580350
rect -736 580294 -680 580350
rect -612 580294 -556 580350
rect -488 580294 -432 580350
rect -860 580170 -804 580226
rect -736 580170 -680 580226
rect -612 580170 -556 580226
rect -488 580170 -432 580226
rect -860 580046 -804 580102
rect -736 580046 -680 580102
rect -612 580046 -556 580102
rect -488 580046 -432 580102
rect -860 579922 -804 579978
rect -736 579922 -680 579978
rect -612 579922 -556 579978
rect -488 579922 -432 579978
rect -860 562294 -804 562350
rect -736 562294 -680 562350
rect -612 562294 -556 562350
rect -488 562294 -432 562350
rect -860 562170 -804 562226
rect -736 562170 -680 562226
rect -612 562170 -556 562226
rect -488 562170 -432 562226
rect -860 562046 -804 562102
rect -736 562046 -680 562102
rect -612 562046 -556 562102
rect -488 562046 -432 562102
rect -860 561922 -804 561978
rect -736 561922 -680 561978
rect -612 561922 -556 561978
rect -488 561922 -432 561978
rect -860 544294 -804 544350
rect -736 544294 -680 544350
rect -612 544294 -556 544350
rect -488 544294 -432 544350
rect -860 544170 -804 544226
rect -736 544170 -680 544226
rect -612 544170 -556 544226
rect -488 544170 -432 544226
rect -860 544046 -804 544102
rect -736 544046 -680 544102
rect -612 544046 -556 544102
rect -488 544046 -432 544102
rect -860 543922 -804 543978
rect -736 543922 -680 543978
rect -612 543922 -556 543978
rect -488 543922 -432 543978
rect -860 526294 -804 526350
rect -736 526294 -680 526350
rect -612 526294 -556 526350
rect -488 526294 -432 526350
rect -860 526170 -804 526226
rect -736 526170 -680 526226
rect -612 526170 -556 526226
rect -488 526170 -432 526226
rect -860 526046 -804 526102
rect -736 526046 -680 526102
rect -612 526046 -556 526102
rect -488 526046 -432 526102
rect -860 525922 -804 525978
rect -736 525922 -680 525978
rect -612 525922 -556 525978
rect -488 525922 -432 525978
rect -860 508294 -804 508350
rect -736 508294 -680 508350
rect -612 508294 -556 508350
rect -488 508294 -432 508350
rect -860 508170 -804 508226
rect -736 508170 -680 508226
rect -612 508170 -556 508226
rect -488 508170 -432 508226
rect -860 508046 -804 508102
rect -736 508046 -680 508102
rect -612 508046 -556 508102
rect -488 508046 -432 508102
rect -860 507922 -804 507978
rect -736 507922 -680 507978
rect -612 507922 -556 507978
rect -488 507922 -432 507978
rect -860 490294 -804 490350
rect -736 490294 -680 490350
rect -612 490294 -556 490350
rect -488 490294 -432 490350
rect -860 490170 -804 490226
rect -736 490170 -680 490226
rect -612 490170 -556 490226
rect -488 490170 -432 490226
rect -860 490046 -804 490102
rect -736 490046 -680 490102
rect -612 490046 -556 490102
rect -488 490046 -432 490102
rect -860 489922 -804 489978
rect -736 489922 -680 489978
rect -612 489922 -556 489978
rect -488 489922 -432 489978
rect -860 472294 -804 472350
rect -736 472294 -680 472350
rect -612 472294 -556 472350
rect -488 472294 -432 472350
rect -860 472170 -804 472226
rect -736 472170 -680 472226
rect -612 472170 -556 472226
rect -488 472170 -432 472226
rect -860 472046 -804 472102
rect -736 472046 -680 472102
rect -612 472046 -556 472102
rect -488 472046 -432 472102
rect -860 471922 -804 471978
rect -736 471922 -680 471978
rect -612 471922 -556 471978
rect -488 471922 -432 471978
rect -860 454294 -804 454350
rect -736 454294 -680 454350
rect -612 454294 -556 454350
rect -488 454294 -432 454350
rect -860 454170 -804 454226
rect -736 454170 -680 454226
rect -612 454170 -556 454226
rect -488 454170 -432 454226
rect -860 454046 -804 454102
rect -736 454046 -680 454102
rect -612 454046 -556 454102
rect -488 454046 -432 454102
rect -860 453922 -804 453978
rect -736 453922 -680 453978
rect -612 453922 -556 453978
rect -488 453922 -432 453978
rect -860 436294 -804 436350
rect -736 436294 -680 436350
rect -612 436294 -556 436350
rect -488 436294 -432 436350
rect -860 436170 -804 436226
rect -736 436170 -680 436226
rect -612 436170 -556 436226
rect -488 436170 -432 436226
rect -860 436046 -804 436102
rect -736 436046 -680 436102
rect -612 436046 -556 436102
rect -488 436046 -432 436102
rect -860 435922 -804 435978
rect -736 435922 -680 435978
rect -612 435922 -556 435978
rect -488 435922 -432 435978
rect -860 418294 -804 418350
rect -736 418294 -680 418350
rect -612 418294 -556 418350
rect -488 418294 -432 418350
rect -860 418170 -804 418226
rect -736 418170 -680 418226
rect -612 418170 -556 418226
rect -488 418170 -432 418226
rect -860 418046 -804 418102
rect -736 418046 -680 418102
rect -612 418046 -556 418102
rect -488 418046 -432 418102
rect -860 417922 -804 417978
rect -736 417922 -680 417978
rect -612 417922 -556 417978
rect -488 417922 -432 417978
rect -860 400294 -804 400350
rect -736 400294 -680 400350
rect -612 400294 -556 400350
rect -488 400294 -432 400350
rect -860 400170 -804 400226
rect -736 400170 -680 400226
rect -612 400170 -556 400226
rect -488 400170 -432 400226
rect -860 400046 -804 400102
rect -736 400046 -680 400102
rect -612 400046 -556 400102
rect -488 400046 -432 400102
rect -860 399922 -804 399978
rect -736 399922 -680 399978
rect -612 399922 -556 399978
rect -488 399922 -432 399978
rect -860 382294 -804 382350
rect -736 382294 -680 382350
rect -612 382294 -556 382350
rect -488 382294 -432 382350
rect -860 382170 -804 382226
rect -736 382170 -680 382226
rect -612 382170 -556 382226
rect -488 382170 -432 382226
rect -860 382046 -804 382102
rect -736 382046 -680 382102
rect -612 382046 -556 382102
rect -488 382046 -432 382102
rect -860 381922 -804 381978
rect -736 381922 -680 381978
rect -612 381922 -556 381978
rect -488 381922 -432 381978
rect -860 364294 -804 364350
rect -736 364294 -680 364350
rect -612 364294 -556 364350
rect -488 364294 -432 364350
rect -860 364170 -804 364226
rect -736 364170 -680 364226
rect -612 364170 -556 364226
rect -488 364170 -432 364226
rect -860 364046 -804 364102
rect -736 364046 -680 364102
rect -612 364046 -556 364102
rect -488 364046 -432 364102
rect -860 363922 -804 363978
rect -736 363922 -680 363978
rect -612 363922 -556 363978
rect -488 363922 -432 363978
rect -860 346294 -804 346350
rect -736 346294 -680 346350
rect -612 346294 -556 346350
rect -488 346294 -432 346350
rect -860 346170 -804 346226
rect -736 346170 -680 346226
rect -612 346170 -556 346226
rect -488 346170 -432 346226
rect -860 346046 -804 346102
rect -736 346046 -680 346102
rect -612 346046 -556 346102
rect -488 346046 -432 346102
rect -860 345922 -804 345978
rect -736 345922 -680 345978
rect -612 345922 -556 345978
rect -488 345922 -432 345978
rect -860 328294 -804 328350
rect -736 328294 -680 328350
rect -612 328294 -556 328350
rect -488 328294 -432 328350
rect -860 328170 -804 328226
rect -736 328170 -680 328226
rect -612 328170 -556 328226
rect -488 328170 -432 328226
rect -860 328046 -804 328102
rect -736 328046 -680 328102
rect -612 328046 -556 328102
rect -488 328046 -432 328102
rect -860 327922 -804 327978
rect -736 327922 -680 327978
rect -612 327922 -556 327978
rect -488 327922 -432 327978
rect -860 310294 -804 310350
rect -736 310294 -680 310350
rect -612 310294 -556 310350
rect -488 310294 -432 310350
rect -860 310170 -804 310226
rect -736 310170 -680 310226
rect -612 310170 -556 310226
rect -488 310170 -432 310226
rect -860 310046 -804 310102
rect -736 310046 -680 310102
rect -612 310046 -556 310102
rect -488 310046 -432 310102
rect -860 309922 -804 309978
rect -736 309922 -680 309978
rect -612 309922 -556 309978
rect -488 309922 -432 309978
rect -860 292294 -804 292350
rect -736 292294 -680 292350
rect -612 292294 -556 292350
rect -488 292294 -432 292350
rect -860 292170 -804 292226
rect -736 292170 -680 292226
rect -612 292170 -556 292226
rect -488 292170 -432 292226
rect -860 292046 -804 292102
rect -736 292046 -680 292102
rect -612 292046 -556 292102
rect -488 292046 -432 292102
rect -860 291922 -804 291978
rect -736 291922 -680 291978
rect -612 291922 -556 291978
rect -488 291922 -432 291978
rect -860 274294 -804 274350
rect -736 274294 -680 274350
rect -612 274294 -556 274350
rect -488 274294 -432 274350
rect -860 274170 -804 274226
rect -736 274170 -680 274226
rect -612 274170 -556 274226
rect -488 274170 -432 274226
rect -860 274046 -804 274102
rect -736 274046 -680 274102
rect -612 274046 -556 274102
rect -488 274046 -432 274102
rect -860 273922 -804 273978
rect -736 273922 -680 273978
rect -612 273922 -556 273978
rect -488 273922 -432 273978
rect -860 256294 -804 256350
rect -736 256294 -680 256350
rect -612 256294 -556 256350
rect -488 256294 -432 256350
rect -860 256170 -804 256226
rect -736 256170 -680 256226
rect -612 256170 -556 256226
rect -488 256170 -432 256226
rect -860 256046 -804 256102
rect -736 256046 -680 256102
rect -612 256046 -556 256102
rect -488 256046 -432 256102
rect -860 255922 -804 255978
rect -736 255922 -680 255978
rect -612 255922 -556 255978
rect -488 255922 -432 255978
rect -860 238294 -804 238350
rect -736 238294 -680 238350
rect -612 238294 -556 238350
rect -488 238294 -432 238350
rect -860 238170 -804 238226
rect -736 238170 -680 238226
rect -612 238170 -556 238226
rect -488 238170 -432 238226
rect -860 238046 -804 238102
rect -736 238046 -680 238102
rect -612 238046 -556 238102
rect -488 238046 -432 238102
rect -860 237922 -804 237978
rect -736 237922 -680 237978
rect -612 237922 -556 237978
rect -488 237922 -432 237978
rect -860 220294 -804 220350
rect -736 220294 -680 220350
rect -612 220294 -556 220350
rect -488 220294 -432 220350
rect -860 220170 -804 220226
rect -736 220170 -680 220226
rect -612 220170 -556 220226
rect -488 220170 -432 220226
rect -860 220046 -804 220102
rect -736 220046 -680 220102
rect -612 220046 -556 220102
rect -488 220046 -432 220102
rect -860 219922 -804 219978
rect -736 219922 -680 219978
rect -612 219922 -556 219978
rect -488 219922 -432 219978
rect -860 202294 -804 202350
rect -736 202294 -680 202350
rect -612 202294 -556 202350
rect -488 202294 -432 202350
rect -860 202170 -804 202226
rect -736 202170 -680 202226
rect -612 202170 -556 202226
rect -488 202170 -432 202226
rect -860 202046 -804 202102
rect -736 202046 -680 202102
rect -612 202046 -556 202102
rect -488 202046 -432 202102
rect -860 201922 -804 201978
rect -736 201922 -680 201978
rect -612 201922 -556 201978
rect -488 201922 -432 201978
rect -860 184294 -804 184350
rect -736 184294 -680 184350
rect -612 184294 -556 184350
rect -488 184294 -432 184350
rect -860 184170 -804 184226
rect -736 184170 -680 184226
rect -612 184170 -556 184226
rect -488 184170 -432 184226
rect -860 184046 -804 184102
rect -736 184046 -680 184102
rect -612 184046 -556 184102
rect -488 184046 -432 184102
rect -860 183922 -804 183978
rect -736 183922 -680 183978
rect -612 183922 -556 183978
rect -488 183922 -432 183978
rect -860 166294 -804 166350
rect -736 166294 -680 166350
rect -612 166294 -556 166350
rect -488 166294 -432 166350
rect -860 166170 -804 166226
rect -736 166170 -680 166226
rect -612 166170 -556 166226
rect -488 166170 -432 166226
rect -860 166046 -804 166102
rect -736 166046 -680 166102
rect -612 166046 -556 166102
rect -488 166046 -432 166102
rect -860 165922 -804 165978
rect -736 165922 -680 165978
rect -612 165922 -556 165978
rect -488 165922 -432 165978
rect -860 148294 -804 148350
rect -736 148294 -680 148350
rect -612 148294 -556 148350
rect -488 148294 -432 148350
rect -860 148170 -804 148226
rect -736 148170 -680 148226
rect -612 148170 -556 148226
rect -488 148170 -432 148226
rect -860 148046 -804 148102
rect -736 148046 -680 148102
rect -612 148046 -556 148102
rect -488 148046 -432 148102
rect -860 147922 -804 147978
rect -736 147922 -680 147978
rect -612 147922 -556 147978
rect -488 147922 -432 147978
rect -860 130294 -804 130350
rect -736 130294 -680 130350
rect -612 130294 -556 130350
rect -488 130294 -432 130350
rect -860 130170 -804 130226
rect -736 130170 -680 130226
rect -612 130170 -556 130226
rect -488 130170 -432 130226
rect -860 130046 -804 130102
rect -736 130046 -680 130102
rect -612 130046 -556 130102
rect -488 130046 -432 130102
rect -860 129922 -804 129978
rect -736 129922 -680 129978
rect -612 129922 -556 129978
rect -488 129922 -432 129978
rect -860 112294 -804 112350
rect -736 112294 -680 112350
rect -612 112294 -556 112350
rect -488 112294 -432 112350
rect -860 112170 -804 112226
rect -736 112170 -680 112226
rect -612 112170 -556 112226
rect -488 112170 -432 112226
rect -860 112046 -804 112102
rect -736 112046 -680 112102
rect -612 112046 -556 112102
rect -488 112046 -432 112102
rect -860 111922 -804 111978
rect -736 111922 -680 111978
rect -612 111922 -556 111978
rect -488 111922 -432 111978
rect -860 94294 -804 94350
rect -736 94294 -680 94350
rect -612 94294 -556 94350
rect -488 94294 -432 94350
rect -860 94170 -804 94226
rect -736 94170 -680 94226
rect -612 94170 -556 94226
rect -488 94170 -432 94226
rect -860 94046 -804 94102
rect -736 94046 -680 94102
rect -612 94046 -556 94102
rect -488 94046 -432 94102
rect -860 93922 -804 93978
rect -736 93922 -680 93978
rect -612 93922 -556 93978
rect -488 93922 -432 93978
rect -860 76294 -804 76350
rect -736 76294 -680 76350
rect -612 76294 -556 76350
rect -488 76294 -432 76350
rect -860 76170 -804 76226
rect -736 76170 -680 76226
rect -612 76170 -556 76226
rect -488 76170 -432 76226
rect -860 76046 -804 76102
rect -736 76046 -680 76102
rect -612 76046 -556 76102
rect -488 76046 -432 76102
rect -860 75922 -804 75978
rect -736 75922 -680 75978
rect -612 75922 -556 75978
rect -488 75922 -432 75978
rect -860 58294 -804 58350
rect -736 58294 -680 58350
rect -612 58294 -556 58350
rect -488 58294 -432 58350
rect -860 58170 -804 58226
rect -736 58170 -680 58226
rect -612 58170 -556 58226
rect -488 58170 -432 58226
rect -860 58046 -804 58102
rect -736 58046 -680 58102
rect -612 58046 -556 58102
rect -488 58046 -432 58102
rect -860 57922 -804 57978
rect -736 57922 -680 57978
rect -612 57922 -556 57978
rect -488 57922 -432 57978
rect -860 40294 -804 40350
rect -736 40294 -680 40350
rect -612 40294 -556 40350
rect -488 40294 -432 40350
rect -860 40170 -804 40226
rect -736 40170 -680 40226
rect -612 40170 -556 40226
rect -488 40170 -432 40226
rect -860 40046 -804 40102
rect -736 40046 -680 40102
rect -612 40046 -556 40102
rect -488 40046 -432 40102
rect -860 39922 -804 39978
rect -736 39922 -680 39978
rect -612 39922 -556 39978
rect -488 39922 -432 39978
rect -860 22294 -804 22350
rect -736 22294 -680 22350
rect -612 22294 -556 22350
rect -488 22294 -432 22350
rect -860 22170 -804 22226
rect -736 22170 -680 22226
rect -612 22170 -556 22226
rect -488 22170 -432 22226
rect -860 22046 -804 22102
rect -736 22046 -680 22102
rect -612 22046 -556 22102
rect -488 22046 -432 22102
rect -860 21922 -804 21978
rect -736 21922 -680 21978
rect -612 21922 -556 21978
rect -488 21922 -432 21978
rect -860 4294 -804 4350
rect -736 4294 -680 4350
rect -612 4294 -556 4350
rect -488 4294 -432 4350
rect -860 4170 -804 4226
rect -736 4170 -680 4226
rect -612 4170 -556 4226
rect -488 4170 -432 4226
rect -860 4046 -804 4102
rect -736 4046 -680 4102
rect -612 4046 -556 4102
rect -488 4046 -432 4102
rect -860 3922 -804 3978
rect -736 3922 -680 3978
rect -612 3922 -556 3978
rect -488 3922 -432 3978
rect -860 -216 -804 -160
rect -736 -216 -680 -160
rect -612 -216 -556 -160
rect -488 -216 -432 -160
rect -860 -340 -804 -284
rect -736 -340 -680 -284
rect -612 -340 -556 -284
rect -488 -340 -432 -284
rect -860 -464 -804 -408
rect -736 -464 -680 -408
rect -612 -464 -556 -408
rect -488 -464 -432 -408
rect -860 -588 -804 -532
rect -736 -588 -680 -532
rect -612 -588 -556 -532
rect -488 -588 -432 -532
rect 3250 597156 3306 597212
rect 3374 597156 3430 597212
rect 3498 597156 3554 597212
rect 3622 597156 3678 597212
rect 3250 597032 3306 597088
rect 3374 597032 3430 597088
rect 3498 597032 3554 597088
rect 3622 597032 3678 597088
rect 3250 596908 3306 596964
rect 3374 596908 3430 596964
rect 3498 596908 3554 596964
rect 3622 596908 3678 596964
rect 3250 596784 3306 596840
rect 3374 596784 3430 596840
rect 3498 596784 3554 596840
rect 3622 596784 3678 596840
rect 3250 580294 3306 580350
rect 3374 580294 3430 580350
rect 3498 580294 3554 580350
rect 3622 580294 3678 580350
rect 3250 580170 3306 580226
rect 3374 580170 3430 580226
rect 3498 580170 3554 580226
rect 3622 580170 3678 580226
rect 3250 580046 3306 580102
rect 3374 580046 3430 580102
rect 3498 580046 3554 580102
rect 3622 580046 3678 580102
rect 3250 579922 3306 579978
rect 3374 579922 3430 579978
rect 3498 579922 3554 579978
rect 3622 579922 3678 579978
rect 3250 562294 3306 562350
rect 3374 562294 3430 562350
rect 3498 562294 3554 562350
rect 3622 562294 3678 562350
rect 3250 562170 3306 562226
rect 3374 562170 3430 562226
rect 3498 562170 3554 562226
rect 3622 562170 3678 562226
rect 3250 562046 3306 562102
rect 3374 562046 3430 562102
rect 3498 562046 3554 562102
rect 3622 562046 3678 562102
rect 3250 561922 3306 561978
rect 3374 561922 3430 561978
rect 3498 561922 3554 561978
rect 3622 561922 3678 561978
rect 3250 544294 3306 544350
rect 3374 544294 3430 544350
rect 3498 544294 3554 544350
rect 3622 544294 3678 544350
rect 3250 544170 3306 544226
rect 3374 544170 3430 544226
rect 3498 544170 3554 544226
rect 3622 544170 3678 544226
rect 3250 544046 3306 544102
rect 3374 544046 3430 544102
rect 3498 544046 3554 544102
rect 3622 544046 3678 544102
rect 3250 543922 3306 543978
rect 3374 543922 3430 543978
rect 3498 543922 3554 543978
rect 3622 543922 3678 543978
rect 3250 526294 3306 526350
rect 3374 526294 3430 526350
rect 3498 526294 3554 526350
rect 3622 526294 3678 526350
rect 3250 526170 3306 526226
rect 3374 526170 3430 526226
rect 3498 526170 3554 526226
rect 3622 526170 3678 526226
rect 3250 526046 3306 526102
rect 3374 526046 3430 526102
rect 3498 526046 3554 526102
rect 3622 526046 3678 526102
rect 3250 525922 3306 525978
rect 3374 525922 3430 525978
rect 3498 525922 3554 525978
rect 3622 525922 3678 525978
rect 3250 508294 3306 508350
rect 3374 508294 3430 508350
rect 3498 508294 3554 508350
rect 3622 508294 3678 508350
rect 3250 508170 3306 508226
rect 3374 508170 3430 508226
rect 3498 508170 3554 508226
rect 3622 508170 3678 508226
rect 3250 508046 3306 508102
rect 3374 508046 3430 508102
rect 3498 508046 3554 508102
rect 3622 508046 3678 508102
rect 3250 507922 3306 507978
rect 3374 507922 3430 507978
rect 3498 507922 3554 507978
rect 3622 507922 3678 507978
rect 3250 490294 3306 490350
rect 3374 490294 3430 490350
rect 3498 490294 3554 490350
rect 3622 490294 3678 490350
rect 3250 490170 3306 490226
rect 3374 490170 3430 490226
rect 3498 490170 3554 490226
rect 3622 490170 3678 490226
rect 3250 490046 3306 490102
rect 3374 490046 3430 490102
rect 3498 490046 3554 490102
rect 3622 490046 3678 490102
rect 3250 489922 3306 489978
rect 3374 489922 3430 489978
rect 3498 489922 3554 489978
rect 3622 489922 3678 489978
rect 3250 472294 3306 472350
rect 3374 472294 3430 472350
rect 3498 472294 3554 472350
rect 3622 472294 3678 472350
rect 3250 472170 3306 472226
rect 3374 472170 3430 472226
rect 3498 472170 3554 472226
rect 3622 472170 3678 472226
rect 3250 472046 3306 472102
rect 3374 472046 3430 472102
rect 3498 472046 3554 472102
rect 3622 472046 3678 472102
rect 3250 471922 3306 471978
rect 3374 471922 3430 471978
rect 3498 471922 3554 471978
rect 3622 471922 3678 471978
rect 3250 454294 3306 454350
rect 3374 454294 3430 454350
rect 3498 454294 3554 454350
rect 3622 454294 3678 454350
rect 3250 454170 3306 454226
rect 3374 454170 3430 454226
rect 3498 454170 3554 454226
rect 3622 454170 3678 454226
rect 3250 454046 3306 454102
rect 3374 454046 3430 454102
rect 3498 454046 3554 454102
rect 3622 454046 3678 454102
rect 3250 453922 3306 453978
rect 3374 453922 3430 453978
rect 3498 453922 3554 453978
rect 3622 453922 3678 453978
rect 3250 436294 3306 436350
rect 3374 436294 3430 436350
rect 3498 436294 3554 436350
rect 3622 436294 3678 436350
rect 3250 436170 3306 436226
rect 3374 436170 3430 436226
rect 3498 436170 3554 436226
rect 3622 436170 3678 436226
rect 3250 436046 3306 436102
rect 3374 436046 3430 436102
rect 3498 436046 3554 436102
rect 3622 436046 3678 436102
rect 3250 435922 3306 435978
rect 3374 435922 3430 435978
rect 3498 435922 3554 435978
rect 3622 435922 3678 435978
rect 3250 418294 3306 418350
rect 3374 418294 3430 418350
rect 3498 418294 3554 418350
rect 3622 418294 3678 418350
rect 3250 418170 3306 418226
rect 3374 418170 3430 418226
rect 3498 418170 3554 418226
rect 3622 418170 3678 418226
rect 3250 418046 3306 418102
rect 3374 418046 3430 418102
rect 3498 418046 3554 418102
rect 3622 418046 3678 418102
rect 3250 417922 3306 417978
rect 3374 417922 3430 417978
rect 3498 417922 3554 417978
rect 3622 417922 3678 417978
rect 3250 400294 3306 400350
rect 3374 400294 3430 400350
rect 3498 400294 3554 400350
rect 3622 400294 3678 400350
rect 3250 400170 3306 400226
rect 3374 400170 3430 400226
rect 3498 400170 3554 400226
rect 3622 400170 3678 400226
rect 3250 400046 3306 400102
rect 3374 400046 3430 400102
rect 3498 400046 3554 400102
rect 3622 400046 3678 400102
rect 3250 399922 3306 399978
rect 3374 399922 3430 399978
rect 3498 399922 3554 399978
rect 3622 399922 3678 399978
rect 3250 382294 3306 382350
rect 3374 382294 3430 382350
rect 3498 382294 3554 382350
rect 3622 382294 3678 382350
rect 3250 382170 3306 382226
rect 3374 382170 3430 382226
rect 3498 382170 3554 382226
rect 3622 382170 3678 382226
rect 3250 382046 3306 382102
rect 3374 382046 3430 382102
rect 3498 382046 3554 382102
rect 3622 382046 3678 382102
rect 3250 381922 3306 381978
rect 3374 381922 3430 381978
rect 3498 381922 3554 381978
rect 3622 381922 3678 381978
rect 3250 364294 3306 364350
rect 3374 364294 3430 364350
rect 3498 364294 3554 364350
rect 3622 364294 3678 364350
rect 3250 364170 3306 364226
rect 3374 364170 3430 364226
rect 3498 364170 3554 364226
rect 3622 364170 3678 364226
rect 3250 364046 3306 364102
rect 3374 364046 3430 364102
rect 3498 364046 3554 364102
rect 3622 364046 3678 364102
rect 3250 363922 3306 363978
rect 3374 363922 3430 363978
rect 3498 363922 3554 363978
rect 3622 363922 3678 363978
rect 3250 346294 3306 346350
rect 3374 346294 3430 346350
rect 3498 346294 3554 346350
rect 3622 346294 3678 346350
rect 3250 346170 3306 346226
rect 3374 346170 3430 346226
rect 3498 346170 3554 346226
rect 3622 346170 3678 346226
rect 3250 346046 3306 346102
rect 3374 346046 3430 346102
rect 3498 346046 3554 346102
rect 3622 346046 3678 346102
rect 3250 345922 3306 345978
rect 3374 345922 3430 345978
rect 3498 345922 3554 345978
rect 3622 345922 3678 345978
rect 3250 328294 3306 328350
rect 3374 328294 3430 328350
rect 3498 328294 3554 328350
rect 3622 328294 3678 328350
rect 3250 328170 3306 328226
rect 3374 328170 3430 328226
rect 3498 328170 3554 328226
rect 3622 328170 3678 328226
rect 3250 328046 3306 328102
rect 3374 328046 3430 328102
rect 3498 328046 3554 328102
rect 3622 328046 3678 328102
rect 3250 327922 3306 327978
rect 3374 327922 3430 327978
rect 3498 327922 3554 327978
rect 3622 327922 3678 327978
rect 3250 310294 3306 310350
rect 3374 310294 3430 310350
rect 3498 310294 3554 310350
rect 3622 310294 3678 310350
rect 3250 310170 3306 310226
rect 3374 310170 3430 310226
rect 3498 310170 3554 310226
rect 3622 310170 3678 310226
rect 3250 310046 3306 310102
rect 3374 310046 3430 310102
rect 3498 310046 3554 310102
rect 3622 310046 3678 310102
rect 3250 309922 3306 309978
rect 3374 309922 3430 309978
rect 3498 309922 3554 309978
rect 3622 309922 3678 309978
rect 3250 292294 3306 292350
rect 3374 292294 3430 292350
rect 3498 292294 3554 292350
rect 3622 292294 3678 292350
rect 3250 292170 3306 292226
rect 3374 292170 3430 292226
rect 3498 292170 3554 292226
rect 3622 292170 3678 292226
rect 3250 292046 3306 292102
rect 3374 292046 3430 292102
rect 3498 292046 3554 292102
rect 3622 292046 3678 292102
rect 3250 291922 3306 291978
rect 3374 291922 3430 291978
rect 3498 291922 3554 291978
rect 3622 291922 3678 291978
rect 3250 274294 3306 274350
rect 3374 274294 3430 274350
rect 3498 274294 3554 274350
rect 3622 274294 3678 274350
rect 3250 274170 3306 274226
rect 3374 274170 3430 274226
rect 3498 274170 3554 274226
rect 3622 274170 3678 274226
rect 3250 274046 3306 274102
rect 3374 274046 3430 274102
rect 3498 274046 3554 274102
rect 3622 274046 3678 274102
rect 3250 273922 3306 273978
rect 3374 273922 3430 273978
rect 3498 273922 3554 273978
rect 3622 273922 3678 273978
rect 3250 256294 3306 256350
rect 3374 256294 3430 256350
rect 3498 256294 3554 256350
rect 3622 256294 3678 256350
rect 3250 256170 3306 256226
rect 3374 256170 3430 256226
rect 3498 256170 3554 256226
rect 3622 256170 3678 256226
rect 3250 256046 3306 256102
rect 3374 256046 3430 256102
rect 3498 256046 3554 256102
rect 3622 256046 3678 256102
rect 3250 255922 3306 255978
rect 3374 255922 3430 255978
rect 3498 255922 3554 255978
rect 3622 255922 3678 255978
rect 3250 238294 3306 238350
rect 3374 238294 3430 238350
rect 3498 238294 3554 238350
rect 3622 238294 3678 238350
rect 3250 238170 3306 238226
rect 3374 238170 3430 238226
rect 3498 238170 3554 238226
rect 3622 238170 3678 238226
rect 3250 238046 3306 238102
rect 3374 238046 3430 238102
rect 3498 238046 3554 238102
rect 3622 238046 3678 238102
rect 3250 237922 3306 237978
rect 3374 237922 3430 237978
rect 3498 237922 3554 237978
rect 3622 237922 3678 237978
rect 3250 220294 3306 220350
rect 3374 220294 3430 220350
rect 3498 220294 3554 220350
rect 3622 220294 3678 220350
rect 3250 220170 3306 220226
rect 3374 220170 3430 220226
rect 3498 220170 3554 220226
rect 3622 220170 3678 220226
rect 3250 220046 3306 220102
rect 3374 220046 3430 220102
rect 3498 220046 3554 220102
rect 3622 220046 3678 220102
rect 3250 219922 3306 219978
rect 3374 219922 3430 219978
rect 3498 219922 3554 219978
rect 3622 219922 3678 219978
rect 3250 202294 3306 202350
rect 3374 202294 3430 202350
rect 3498 202294 3554 202350
rect 3622 202294 3678 202350
rect 3250 202170 3306 202226
rect 3374 202170 3430 202226
rect 3498 202170 3554 202226
rect 3622 202170 3678 202226
rect 3250 202046 3306 202102
rect 3374 202046 3430 202102
rect 3498 202046 3554 202102
rect 3622 202046 3678 202102
rect 3250 201922 3306 201978
rect 3374 201922 3430 201978
rect 3498 201922 3554 201978
rect 3622 201922 3678 201978
rect 3250 184294 3306 184350
rect 3374 184294 3430 184350
rect 3498 184294 3554 184350
rect 3622 184294 3678 184350
rect 3250 184170 3306 184226
rect 3374 184170 3430 184226
rect 3498 184170 3554 184226
rect 3622 184170 3678 184226
rect 3250 184046 3306 184102
rect 3374 184046 3430 184102
rect 3498 184046 3554 184102
rect 3622 184046 3678 184102
rect 3250 183922 3306 183978
rect 3374 183922 3430 183978
rect 3498 183922 3554 183978
rect 3622 183922 3678 183978
rect 3250 166294 3306 166350
rect 3374 166294 3430 166350
rect 3498 166294 3554 166350
rect 3622 166294 3678 166350
rect 3250 166170 3306 166226
rect 3374 166170 3430 166226
rect 3498 166170 3554 166226
rect 3622 166170 3678 166226
rect 3250 166046 3306 166102
rect 3374 166046 3430 166102
rect 3498 166046 3554 166102
rect 3622 166046 3678 166102
rect 3250 165922 3306 165978
rect 3374 165922 3430 165978
rect 3498 165922 3554 165978
rect 3622 165922 3678 165978
rect 3250 148294 3306 148350
rect 3374 148294 3430 148350
rect 3498 148294 3554 148350
rect 3622 148294 3678 148350
rect 3250 148170 3306 148226
rect 3374 148170 3430 148226
rect 3498 148170 3554 148226
rect 3622 148170 3678 148226
rect 3250 148046 3306 148102
rect 3374 148046 3430 148102
rect 3498 148046 3554 148102
rect 3622 148046 3678 148102
rect 3250 147922 3306 147978
rect 3374 147922 3430 147978
rect 3498 147922 3554 147978
rect 3622 147922 3678 147978
rect 3250 130294 3306 130350
rect 3374 130294 3430 130350
rect 3498 130294 3554 130350
rect 3622 130294 3678 130350
rect 3250 130170 3306 130226
rect 3374 130170 3430 130226
rect 3498 130170 3554 130226
rect 3622 130170 3678 130226
rect 3250 130046 3306 130102
rect 3374 130046 3430 130102
rect 3498 130046 3554 130102
rect 3622 130046 3678 130102
rect 3250 129922 3306 129978
rect 3374 129922 3430 129978
rect 3498 129922 3554 129978
rect 3622 129922 3678 129978
rect 3250 112294 3306 112350
rect 3374 112294 3430 112350
rect 3498 112294 3554 112350
rect 3622 112294 3678 112350
rect 3250 112170 3306 112226
rect 3374 112170 3430 112226
rect 3498 112170 3554 112226
rect 3622 112170 3678 112226
rect 3250 112046 3306 112102
rect 3374 112046 3430 112102
rect 3498 112046 3554 112102
rect 3622 112046 3678 112102
rect 3250 111922 3306 111978
rect 3374 111922 3430 111978
rect 3498 111922 3554 111978
rect 3622 111922 3678 111978
rect 3250 94294 3306 94350
rect 3374 94294 3430 94350
rect 3498 94294 3554 94350
rect 3622 94294 3678 94350
rect 3250 94170 3306 94226
rect 3374 94170 3430 94226
rect 3498 94170 3554 94226
rect 3622 94170 3678 94226
rect 3250 94046 3306 94102
rect 3374 94046 3430 94102
rect 3498 94046 3554 94102
rect 3622 94046 3678 94102
rect 3250 93922 3306 93978
rect 3374 93922 3430 93978
rect 3498 93922 3554 93978
rect 3622 93922 3678 93978
rect 3250 76294 3306 76350
rect 3374 76294 3430 76350
rect 3498 76294 3554 76350
rect 3622 76294 3678 76350
rect 3250 76170 3306 76226
rect 3374 76170 3430 76226
rect 3498 76170 3554 76226
rect 3622 76170 3678 76226
rect 3250 76046 3306 76102
rect 3374 76046 3430 76102
rect 3498 76046 3554 76102
rect 3622 76046 3678 76102
rect 3250 75922 3306 75978
rect 3374 75922 3430 75978
rect 3498 75922 3554 75978
rect 3622 75922 3678 75978
rect 3250 58294 3306 58350
rect 3374 58294 3430 58350
rect 3498 58294 3554 58350
rect 3622 58294 3678 58350
rect 3250 58170 3306 58226
rect 3374 58170 3430 58226
rect 3498 58170 3554 58226
rect 3622 58170 3678 58226
rect 3250 58046 3306 58102
rect 3374 58046 3430 58102
rect 3498 58046 3554 58102
rect 3622 58046 3678 58102
rect 3250 57922 3306 57978
rect 3374 57922 3430 57978
rect 3498 57922 3554 57978
rect 3622 57922 3678 57978
rect 3250 40294 3306 40350
rect 3374 40294 3430 40350
rect 3498 40294 3554 40350
rect 3622 40294 3678 40350
rect 3250 40170 3306 40226
rect 3374 40170 3430 40226
rect 3498 40170 3554 40226
rect 3622 40170 3678 40226
rect 3250 40046 3306 40102
rect 3374 40046 3430 40102
rect 3498 40046 3554 40102
rect 3622 40046 3678 40102
rect 3250 39922 3306 39978
rect 3374 39922 3430 39978
rect 3498 39922 3554 39978
rect 3622 39922 3678 39978
rect 3250 22294 3306 22350
rect 3374 22294 3430 22350
rect 3498 22294 3554 22350
rect 3622 22294 3678 22350
rect 3250 22170 3306 22226
rect 3374 22170 3430 22226
rect 3498 22170 3554 22226
rect 3622 22170 3678 22226
rect 3250 22046 3306 22102
rect 3374 22046 3430 22102
rect 3498 22046 3554 22102
rect 3622 22046 3678 22102
rect 3250 21922 3306 21978
rect 3374 21922 3430 21978
rect 3498 21922 3554 21978
rect 3622 21922 3678 21978
rect 3250 4294 3306 4350
rect 3374 4294 3430 4350
rect 3498 4294 3554 4350
rect 3622 4294 3678 4350
rect 3250 4170 3306 4226
rect 3374 4170 3430 4226
rect 3498 4170 3554 4226
rect 3622 4170 3678 4226
rect 3250 4046 3306 4102
rect 3374 4046 3430 4102
rect 3498 4046 3554 4102
rect 3622 4046 3678 4102
rect 3250 3922 3306 3978
rect 3374 3922 3430 3978
rect 3498 3922 3554 3978
rect 3622 3922 3678 3978
rect 3250 -216 3306 -160
rect 3374 -216 3430 -160
rect 3498 -216 3554 -160
rect 3622 -216 3678 -160
rect 3250 -340 3306 -284
rect 3374 -340 3430 -284
rect 3498 -340 3554 -284
rect 3622 -340 3678 -284
rect 3250 -464 3306 -408
rect 3374 -464 3430 -408
rect 3498 -464 3554 -408
rect 3622 -464 3678 -408
rect 3250 -588 3306 -532
rect 3374 -588 3430 -532
rect 3498 -588 3554 -532
rect 3622 -588 3678 -532
rect -1820 -1176 -1764 -1120
rect -1696 -1176 -1640 -1120
rect -1572 -1176 -1516 -1120
rect -1448 -1176 -1392 -1120
rect -1820 -1300 -1764 -1244
rect -1696 -1300 -1640 -1244
rect -1572 -1300 -1516 -1244
rect -1448 -1300 -1392 -1244
rect -1820 -1424 -1764 -1368
rect -1696 -1424 -1640 -1368
rect -1572 -1424 -1516 -1368
rect -1448 -1424 -1392 -1368
rect -1820 -1548 -1764 -1492
rect -1696 -1548 -1640 -1492
rect -1572 -1548 -1516 -1492
rect -1448 -1548 -1392 -1492
rect 6970 598116 7026 598172
rect 7094 598116 7150 598172
rect 7218 598116 7274 598172
rect 7342 598116 7398 598172
rect 6970 597992 7026 598048
rect 7094 597992 7150 598048
rect 7218 597992 7274 598048
rect 7342 597992 7398 598048
rect 6970 597868 7026 597924
rect 7094 597868 7150 597924
rect 7218 597868 7274 597924
rect 7342 597868 7398 597924
rect 6970 597744 7026 597800
rect 7094 597744 7150 597800
rect 7218 597744 7274 597800
rect 7342 597744 7398 597800
rect 6970 586294 7026 586350
rect 7094 586294 7150 586350
rect 7218 586294 7274 586350
rect 7342 586294 7398 586350
rect 6970 586170 7026 586226
rect 7094 586170 7150 586226
rect 7218 586170 7274 586226
rect 7342 586170 7398 586226
rect 6970 586046 7026 586102
rect 7094 586046 7150 586102
rect 7218 586046 7274 586102
rect 7342 586046 7398 586102
rect 6970 585922 7026 585978
rect 7094 585922 7150 585978
rect 7218 585922 7274 585978
rect 7342 585922 7398 585978
rect 6970 568294 7026 568350
rect 7094 568294 7150 568350
rect 7218 568294 7274 568350
rect 7342 568294 7398 568350
rect 6970 568170 7026 568226
rect 7094 568170 7150 568226
rect 7218 568170 7274 568226
rect 7342 568170 7398 568226
rect 6970 568046 7026 568102
rect 7094 568046 7150 568102
rect 7218 568046 7274 568102
rect 7342 568046 7398 568102
rect 6970 567922 7026 567978
rect 7094 567922 7150 567978
rect 7218 567922 7274 567978
rect 7342 567922 7398 567978
rect 6970 550294 7026 550350
rect 7094 550294 7150 550350
rect 7218 550294 7274 550350
rect 7342 550294 7398 550350
rect 6970 550170 7026 550226
rect 7094 550170 7150 550226
rect 7218 550170 7274 550226
rect 7342 550170 7398 550226
rect 6970 550046 7026 550102
rect 7094 550046 7150 550102
rect 7218 550046 7274 550102
rect 7342 550046 7398 550102
rect 6970 549922 7026 549978
rect 7094 549922 7150 549978
rect 7218 549922 7274 549978
rect 7342 549922 7398 549978
rect 6970 532294 7026 532350
rect 7094 532294 7150 532350
rect 7218 532294 7274 532350
rect 7342 532294 7398 532350
rect 6970 532170 7026 532226
rect 7094 532170 7150 532226
rect 7218 532170 7274 532226
rect 7342 532170 7398 532226
rect 6970 532046 7026 532102
rect 7094 532046 7150 532102
rect 7218 532046 7274 532102
rect 7342 532046 7398 532102
rect 6970 531922 7026 531978
rect 7094 531922 7150 531978
rect 7218 531922 7274 531978
rect 7342 531922 7398 531978
rect 6970 514294 7026 514350
rect 7094 514294 7150 514350
rect 7218 514294 7274 514350
rect 7342 514294 7398 514350
rect 6970 514170 7026 514226
rect 7094 514170 7150 514226
rect 7218 514170 7274 514226
rect 7342 514170 7398 514226
rect 6970 514046 7026 514102
rect 7094 514046 7150 514102
rect 7218 514046 7274 514102
rect 7342 514046 7398 514102
rect 6970 513922 7026 513978
rect 7094 513922 7150 513978
rect 7218 513922 7274 513978
rect 7342 513922 7398 513978
rect 6970 496294 7026 496350
rect 7094 496294 7150 496350
rect 7218 496294 7274 496350
rect 7342 496294 7398 496350
rect 6970 496170 7026 496226
rect 7094 496170 7150 496226
rect 7218 496170 7274 496226
rect 7342 496170 7398 496226
rect 6970 496046 7026 496102
rect 7094 496046 7150 496102
rect 7218 496046 7274 496102
rect 7342 496046 7398 496102
rect 6970 495922 7026 495978
rect 7094 495922 7150 495978
rect 7218 495922 7274 495978
rect 7342 495922 7398 495978
rect 6970 478294 7026 478350
rect 7094 478294 7150 478350
rect 7218 478294 7274 478350
rect 7342 478294 7398 478350
rect 6970 478170 7026 478226
rect 7094 478170 7150 478226
rect 7218 478170 7274 478226
rect 7342 478170 7398 478226
rect 6970 478046 7026 478102
rect 7094 478046 7150 478102
rect 7218 478046 7274 478102
rect 7342 478046 7398 478102
rect 6970 477922 7026 477978
rect 7094 477922 7150 477978
rect 7218 477922 7274 477978
rect 7342 477922 7398 477978
rect 6970 460294 7026 460350
rect 7094 460294 7150 460350
rect 7218 460294 7274 460350
rect 7342 460294 7398 460350
rect 6970 460170 7026 460226
rect 7094 460170 7150 460226
rect 7218 460170 7274 460226
rect 7342 460170 7398 460226
rect 6970 460046 7026 460102
rect 7094 460046 7150 460102
rect 7218 460046 7274 460102
rect 7342 460046 7398 460102
rect 6970 459922 7026 459978
rect 7094 459922 7150 459978
rect 7218 459922 7274 459978
rect 7342 459922 7398 459978
rect 6970 442294 7026 442350
rect 7094 442294 7150 442350
rect 7218 442294 7274 442350
rect 7342 442294 7398 442350
rect 6970 442170 7026 442226
rect 7094 442170 7150 442226
rect 7218 442170 7274 442226
rect 7342 442170 7398 442226
rect 6970 442046 7026 442102
rect 7094 442046 7150 442102
rect 7218 442046 7274 442102
rect 7342 442046 7398 442102
rect 6970 441922 7026 441978
rect 7094 441922 7150 441978
rect 7218 441922 7274 441978
rect 7342 441922 7398 441978
rect 6970 424294 7026 424350
rect 7094 424294 7150 424350
rect 7218 424294 7274 424350
rect 7342 424294 7398 424350
rect 6970 424170 7026 424226
rect 7094 424170 7150 424226
rect 7218 424170 7274 424226
rect 7342 424170 7398 424226
rect 6970 424046 7026 424102
rect 7094 424046 7150 424102
rect 7218 424046 7274 424102
rect 7342 424046 7398 424102
rect 6970 423922 7026 423978
rect 7094 423922 7150 423978
rect 7218 423922 7274 423978
rect 7342 423922 7398 423978
rect 6970 406294 7026 406350
rect 7094 406294 7150 406350
rect 7218 406294 7274 406350
rect 7342 406294 7398 406350
rect 6970 406170 7026 406226
rect 7094 406170 7150 406226
rect 7218 406170 7274 406226
rect 7342 406170 7398 406226
rect 6970 406046 7026 406102
rect 7094 406046 7150 406102
rect 7218 406046 7274 406102
rect 7342 406046 7398 406102
rect 6970 405922 7026 405978
rect 7094 405922 7150 405978
rect 7218 405922 7274 405978
rect 7342 405922 7398 405978
rect 6970 388294 7026 388350
rect 7094 388294 7150 388350
rect 7218 388294 7274 388350
rect 7342 388294 7398 388350
rect 6970 388170 7026 388226
rect 7094 388170 7150 388226
rect 7218 388170 7274 388226
rect 7342 388170 7398 388226
rect 6970 388046 7026 388102
rect 7094 388046 7150 388102
rect 7218 388046 7274 388102
rect 7342 388046 7398 388102
rect 6970 387922 7026 387978
rect 7094 387922 7150 387978
rect 7218 387922 7274 387978
rect 7342 387922 7398 387978
rect 6970 370294 7026 370350
rect 7094 370294 7150 370350
rect 7218 370294 7274 370350
rect 7342 370294 7398 370350
rect 6970 370170 7026 370226
rect 7094 370170 7150 370226
rect 7218 370170 7274 370226
rect 7342 370170 7398 370226
rect 6970 370046 7026 370102
rect 7094 370046 7150 370102
rect 7218 370046 7274 370102
rect 7342 370046 7398 370102
rect 6970 369922 7026 369978
rect 7094 369922 7150 369978
rect 7218 369922 7274 369978
rect 7342 369922 7398 369978
rect 6970 352294 7026 352350
rect 7094 352294 7150 352350
rect 7218 352294 7274 352350
rect 7342 352294 7398 352350
rect 6970 352170 7026 352226
rect 7094 352170 7150 352226
rect 7218 352170 7274 352226
rect 7342 352170 7398 352226
rect 6970 352046 7026 352102
rect 7094 352046 7150 352102
rect 7218 352046 7274 352102
rect 7342 352046 7398 352102
rect 6970 351922 7026 351978
rect 7094 351922 7150 351978
rect 7218 351922 7274 351978
rect 7342 351922 7398 351978
rect 6970 334294 7026 334350
rect 7094 334294 7150 334350
rect 7218 334294 7274 334350
rect 7342 334294 7398 334350
rect 6970 334170 7026 334226
rect 7094 334170 7150 334226
rect 7218 334170 7274 334226
rect 7342 334170 7398 334226
rect 6970 334046 7026 334102
rect 7094 334046 7150 334102
rect 7218 334046 7274 334102
rect 7342 334046 7398 334102
rect 6970 333922 7026 333978
rect 7094 333922 7150 333978
rect 7218 333922 7274 333978
rect 7342 333922 7398 333978
rect 6970 316294 7026 316350
rect 7094 316294 7150 316350
rect 7218 316294 7274 316350
rect 7342 316294 7398 316350
rect 6970 316170 7026 316226
rect 7094 316170 7150 316226
rect 7218 316170 7274 316226
rect 7342 316170 7398 316226
rect 6970 316046 7026 316102
rect 7094 316046 7150 316102
rect 7218 316046 7274 316102
rect 7342 316046 7398 316102
rect 6970 315922 7026 315978
rect 7094 315922 7150 315978
rect 7218 315922 7274 315978
rect 7342 315922 7398 315978
rect 6970 298294 7026 298350
rect 7094 298294 7150 298350
rect 7218 298294 7274 298350
rect 7342 298294 7398 298350
rect 6970 298170 7026 298226
rect 7094 298170 7150 298226
rect 7218 298170 7274 298226
rect 7342 298170 7398 298226
rect 6970 298046 7026 298102
rect 7094 298046 7150 298102
rect 7218 298046 7274 298102
rect 7342 298046 7398 298102
rect 6970 297922 7026 297978
rect 7094 297922 7150 297978
rect 7218 297922 7274 297978
rect 7342 297922 7398 297978
rect 6970 280294 7026 280350
rect 7094 280294 7150 280350
rect 7218 280294 7274 280350
rect 7342 280294 7398 280350
rect 6970 280170 7026 280226
rect 7094 280170 7150 280226
rect 7218 280170 7274 280226
rect 7342 280170 7398 280226
rect 6970 280046 7026 280102
rect 7094 280046 7150 280102
rect 7218 280046 7274 280102
rect 7342 280046 7398 280102
rect 6970 279922 7026 279978
rect 7094 279922 7150 279978
rect 7218 279922 7274 279978
rect 7342 279922 7398 279978
rect 6970 262294 7026 262350
rect 7094 262294 7150 262350
rect 7218 262294 7274 262350
rect 7342 262294 7398 262350
rect 6970 262170 7026 262226
rect 7094 262170 7150 262226
rect 7218 262170 7274 262226
rect 7342 262170 7398 262226
rect 6970 262046 7026 262102
rect 7094 262046 7150 262102
rect 7218 262046 7274 262102
rect 7342 262046 7398 262102
rect 6970 261922 7026 261978
rect 7094 261922 7150 261978
rect 7218 261922 7274 261978
rect 7342 261922 7398 261978
rect 6970 244294 7026 244350
rect 7094 244294 7150 244350
rect 7218 244294 7274 244350
rect 7342 244294 7398 244350
rect 6970 244170 7026 244226
rect 7094 244170 7150 244226
rect 7218 244170 7274 244226
rect 7342 244170 7398 244226
rect 6970 244046 7026 244102
rect 7094 244046 7150 244102
rect 7218 244046 7274 244102
rect 7342 244046 7398 244102
rect 6970 243922 7026 243978
rect 7094 243922 7150 243978
rect 7218 243922 7274 243978
rect 7342 243922 7398 243978
rect 6970 226294 7026 226350
rect 7094 226294 7150 226350
rect 7218 226294 7274 226350
rect 7342 226294 7398 226350
rect 6970 226170 7026 226226
rect 7094 226170 7150 226226
rect 7218 226170 7274 226226
rect 7342 226170 7398 226226
rect 6970 226046 7026 226102
rect 7094 226046 7150 226102
rect 7218 226046 7274 226102
rect 7342 226046 7398 226102
rect 6970 225922 7026 225978
rect 7094 225922 7150 225978
rect 7218 225922 7274 225978
rect 7342 225922 7398 225978
rect 6970 208294 7026 208350
rect 7094 208294 7150 208350
rect 7218 208294 7274 208350
rect 7342 208294 7398 208350
rect 6970 208170 7026 208226
rect 7094 208170 7150 208226
rect 7218 208170 7274 208226
rect 7342 208170 7398 208226
rect 6970 208046 7026 208102
rect 7094 208046 7150 208102
rect 7218 208046 7274 208102
rect 7342 208046 7398 208102
rect 6970 207922 7026 207978
rect 7094 207922 7150 207978
rect 7218 207922 7274 207978
rect 7342 207922 7398 207978
rect 6970 190294 7026 190350
rect 7094 190294 7150 190350
rect 7218 190294 7274 190350
rect 7342 190294 7398 190350
rect 6970 190170 7026 190226
rect 7094 190170 7150 190226
rect 7218 190170 7274 190226
rect 7342 190170 7398 190226
rect 6970 190046 7026 190102
rect 7094 190046 7150 190102
rect 7218 190046 7274 190102
rect 7342 190046 7398 190102
rect 6970 189922 7026 189978
rect 7094 189922 7150 189978
rect 7218 189922 7274 189978
rect 7342 189922 7398 189978
rect 6970 172294 7026 172350
rect 7094 172294 7150 172350
rect 7218 172294 7274 172350
rect 7342 172294 7398 172350
rect 6970 172170 7026 172226
rect 7094 172170 7150 172226
rect 7218 172170 7274 172226
rect 7342 172170 7398 172226
rect 6970 172046 7026 172102
rect 7094 172046 7150 172102
rect 7218 172046 7274 172102
rect 7342 172046 7398 172102
rect 6970 171922 7026 171978
rect 7094 171922 7150 171978
rect 7218 171922 7274 171978
rect 7342 171922 7398 171978
rect 6970 154294 7026 154350
rect 7094 154294 7150 154350
rect 7218 154294 7274 154350
rect 7342 154294 7398 154350
rect 6970 154170 7026 154226
rect 7094 154170 7150 154226
rect 7218 154170 7274 154226
rect 7342 154170 7398 154226
rect 6970 154046 7026 154102
rect 7094 154046 7150 154102
rect 7218 154046 7274 154102
rect 7342 154046 7398 154102
rect 6970 153922 7026 153978
rect 7094 153922 7150 153978
rect 7218 153922 7274 153978
rect 7342 153922 7398 153978
rect 6970 136294 7026 136350
rect 7094 136294 7150 136350
rect 7218 136294 7274 136350
rect 7342 136294 7398 136350
rect 6970 136170 7026 136226
rect 7094 136170 7150 136226
rect 7218 136170 7274 136226
rect 7342 136170 7398 136226
rect 6970 136046 7026 136102
rect 7094 136046 7150 136102
rect 7218 136046 7274 136102
rect 7342 136046 7398 136102
rect 6970 135922 7026 135978
rect 7094 135922 7150 135978
rect 7218 135922 7274 135978
rect 7342 135922 7398 135978
rect 6970 118294 7026 118350
rect 7094 118294 7150 118350
rect 7218 118294 7274 118350
rect 7342 118294 7398 118350
rect 6970 118170 7026 118226
rect 7094 118170 7150 118226
rect 7218 118170 7274 118226
rect 7342 118170 7398 118226
rect 6970 118046 7026 118102
rect 7094 118046 7150 118102
rect 7218 118046 7274 118102
rect 7342 118046 7398 118102
rect 6970 117922 7026 117978
rect 7094 117922 7150 117978
rect 7218 117922 7274 117978
rect 7342 117922 7398 117978
rect 6970 100294 7026 100350
rect 7094 100294 7150 100350
rect 7218 100294 7274 100350
rect 7342 100294 7398 100350
rect 6970 100170 7026 100226
rect 7094 100170 7150 100226
rect 7218 100170 7274 100226
rect 7342 100170 7398 100226
rect 6970 100046 7026 100102
rect 7094 100046 7150 100102
rect 7218 100046 7274 100102
rect 7342 100046 7398 100102
rect 6970 99922 7026 99978
rect 7094 99922 7150 99978
rect 7218 99922 7274 99978
rect 7342 99922 7398 99978
rect 6970 82294 7026 82350
rect 7094 82294 7150 82350
rect 7218 82294 7274 82350
rect 7342 82294 7398 82350
rect 6970 82170 7026 82226
rect 7094 82170 7150 82226
rect 7218 82170 7274 82226
rect 7342 82170 7398 82226
rect 6970 82046 7026 82102
rect 7094 82046 7150 82102
rect 7218 82046 7274 82102
rect 7342 82046 7398 82102
rect 6970 81922 7026 81978
rect 7094 81922 7150 81978
rect 7218 81922 7274 81978
rect 7342 81922 7398 81978
rect 6970 64294 7026 64350
rect 7094 64294 7150 64350
rect 7218 64294 7274 64350
rect 7342 64294 7398 64350
rect 6970 64170 7026 64226
rect 7094 64170 7150 64226
rect 7218 64170 7274 64226
rect 7342 64170 7398 64226
rect 6970 64046 7026 64102
rect 7094 64046 7150 64102
rect 7218 64046 7274 64102
rect 7342 64046 7398 64102
rect 6970 63922 7026 63978
rect 7094 63922 7150 63978
rect 7218 63922 7274 63978
rect 7342 63922 7398 63978
rect 6970 46294 7026 46350
rect 7094 46294 7150 46350
rect 7218 46294 7274 46350
rect 7342 46294 7398 46350
rect 6970 46170 7026 46226
rect 7094 46170 7150 46226
rect 7218 46170 7274 46226
rect 7342 46170 7398 46226
rect 6970 46046 7026 46102
rect 7094 46046 7150 46102
rect 7218 46046 7274 46102
rect 7342 46046 7398 46102
rect 6970 45922 7026 45978
rect 7094 45922 7150 45978
rect 7218 45922 7274 45978
rect 7342 45922 7398 45978
rect 6970 28294 7026 28350
rect 7094 28294 7150 28350
rect 7218 28294 7274 28350
rect 7342 28294 7398 28350
rect 6970 28170 7026 28226
rect 7094 28170 7150 28226
rect 7218 28170 7274 28226
rect 7342 28170 7398 28226
rect 6970 28046 7026 28102
rect 7094 28046 7150 28102
rect 7218 28046 7274 28102
rect 7342 28046 7398 28102
rect 6970 27922 7026 27978
rect 7094 27922 7150 27978
rect 7218 27922 7274 27978
rect 7342 27922 7398 27978
rect 6970 10294 7026 10350
rect 7094 10294 7150 10350
rect 7218 10294 7274 10350
rect 7342 10294 7398 10350
rect 6970 10170 7026 10226
rect 7094 10170 7150 10226
rect 7218 10170 7274 10226
rect 7342 10170 7398 10226
rect 6970 10046 7026 10102
rect 7094 10046 7150 10102
rect 7218 10046 7274 10102
rect 7342 10046 7398 10102
rect 6970 9922 7026 9978
rect 7094 9922 7150 9978
rect 7218 9922 7274 9978
rect 7342 9922 7398 9978
rect 6970 -1176 7026 -1120
rect 7094 -1176 7150 -1120
rect 7218 -1176 7274 -1120
rect 7342 -1176 7398 -1120
rect 6970 -1300 7026 -1244
rect 7094 -1300 7150 -1244
rect 7218 -1300 7274 -1244
rect 7342 -1300 7398 -1244
rect 6970 -1424 7026 -1368
rect 7094 -1424 7150 -1368
rect 7218 -1424 7274 -1368
rect 7342 -1424 7398 -1368
rect 6970 -1548 7026 -1492
rect 7094 -1548 7150 -1492
rect 7218 -1548 7274 -1492
rect 7342 -1548 7398 -1492
rect 21250 597156 21306 597212
rect 21374 597156 21430 597212
rect 21498 597156 21554 597212
rect 21622 597156 21678 597212
rect 21250 597032 21306 597088
rect 21374 597032 21430 597088
rect 21498 597032 21554 597088
rect 21622 597032 21678 597088
rect 21250 596908 21306 596964
rect 21374 596908 21430 596964
rect 21498 596908 21554 596964
rect 21622 596908 21678 596964
rect 21250 596784 21306 596840
rect 21374 596784 21430 596840
rect 21498 596784 21554 596840
rect 21622 596784 21678 596840
rect 21250 580294 21306 580350
rect 21374 580294 21430 580350
rect 21498 580294 21554 580350
rect 21622 580294 21678 580350
rect 21250 580170 21306 580226
rect 21374 580170 21430 580226
rect 21498 580170 21554 580226
rect 21622 580170 21678 580226
rect 21250 580046 21306 580102
rect 21374 580046 21430 580102
rect 21498 580046 21554 580102
rect 21622 580046 21678 580102
rect 21250 579922 21306 579978
rect 21374 579922 21430 579978
rect 21498 579922 21554 579978
rect 21622 579922 21678 579978
rect 21250 562294 21306 562350
rect 21374 562294 21430 562350
rect 21498 562294 21554 562350
rect 21622 562294 21678 562350
rect 21250 562170 21306 562226
rect 21374 562170 21430 562226
rect 21498 562170 21554 562226
rect 21622 562170 21678 562226
rect 21250 562046 21306 562102
rect 21374 562046 21430 562102
rect 21498 562046 21554 562102
rect 21622 562046 21678 562102
rect 21250 561922 21306 561978
rect 21374 561922 21430 561978
rect 21498 561922 21554 561978
rect 21622 561922 21678 561978
rect 21250 544294 21306 544350
rect 21374 544294 21430 544350
rect 21498 544294 21554 544350
rect 21622 544294 21678 544350
rect 21250 544170 21306 544226
rect 21374 544170 21430 544226
rect 21498 544170 21554 544226
rect 21622 544170 21678 544226
rect 21250 544046 21306 544102
rect 21374 544046 21430 544102
rect 21498 544046 21554 544102
rect 21622 544046 21678 544102
rect 21250 543922 21306 543978
rect 21374 543922 21430 543978
rect 21498 543922 21554 543978
rect 21622 543922 21678 543978
rect 21250 526294 21306 526350
rect 21374 526294 21430 526350
rect 21498 526294 21554 526350
rect 21622 526294 21678 526350
rect 21250 526170 21306 526226
rect 21374 526170 21430 526226
rect 21498 526170 21554 526226
rect 21622 526170 21678 526226
rect 21250 526046 21306 526102
rect 21374 526046 21430 526102
rect 21498 526046 21554 526102
rect 21622 526046 21678 526102
rect 21250 525922 21306 525978
rect 21374 525922 21430 525978
rect 21498 525922 21554 525978
rect 21622 525922 21678 525978
rect 21250 508294 21306 508350
rect 21374 508294 21430 508350
rect 21498 508294 21554 508350
rect 21622 508294 21678 508350
rect 21250 508170 21306 508226
rect 21374 508170 21430 508226
rect 21498 508170 21554 508226
rect 21622 508170 21678 508226
rect 21250 508046 21306 508102
rect 21374 508046 21430 508102
rect 21498 508046 21554 508102
rect 21622 508046 21678 508102
rect 21250 507922 21306 507978
rect 21374 507922 21430 507978
rect 21498 507922 21554 507978
rect 21622 507922 21678 507978
rect 21250 490294 21306 490350
rect 21374 490294 21430 490350
rect 21498 490294 21554 490350
rect 21622 490294 21678 490350
rect 21250 490170 21306 490226
rect 21374 490170 21430 490226
rect 21498 490170 21554 490226
rect 21622 490170 21678 490226
rect 21250 490046 21306 490102
rect 21374 490046 21430 490102
rect 21498 490046 21554 490102
rect 21622 490046 21678 490102
rect 21250 489922 21306 489978
rect 21374 489922 21430 489978
rect 21498 489922 21554 489978
rect 21622 489922 21678 489978
rect 21250 472294 21306 472350
rect 21374 472294 21430 472350
rect 21498 472294 21554 472350
rect 21622 472294 21678 472350
rect 21250 472170 21306 472226
rect 21374 472170 21430 472226
rect 21498 472170 21554 472226
rect 21622 472170 21678 472226
rect 21250 472046 21306 472102
rect 21374 472046 21430 472102
rect 21498 472046 21554 472102
rect 21622 472046 21678 472102
rect 21250 471922 21306 471978
rect 21374 471922 21430 471978
rect 21498 471922 21554 471978
rect 21622 471922 21678 471978
rect 21250 454294 21306 454350
rect 21374 454294 21430 454350
rect 21498 454294 21554 454350
rect 21622 454294 21678 454350
rect 21250 454170 21306 454226
rect 21374 454170 21430 454226
rect 21498 454170 21554 454226
rect 21622 454170 21678 454226
rect 21250 454046 21306 454102
rect 21374 454046 21430 454102
rect 21498 454046 21554 454102
rect 21622 454046 21678 454102
rect 21250 453922 21306 453978
rect 21374 453922 21430 453978
rect 21498 453922 21554 453978
rect 21622 453922 21678 453978
rect 21250 436294 21306 436350
rect 21374 436294 21430 436350
rect 21498 436294 21554 436350
rect 21622 436294 21678 436350
rect 21250 436170 21306 436226
rect 21374 436170 21430 436226
rect 21498 436170 21554 436226
rect 21622 436170 21678 436226
rect 21250 436046 21306 436102
rect 21374 436046 21430 436102
rect 21498 436046 21554 436102
rect 21622 436046 21678 436102
rect 21250 435922 21306 435978
rect 21374 435922 21430 435978
rect 21498 435922 21554 435978
rect 21622 435922 21678 435978
rect 21250 418294 21306 418350
rect 21374 418294 21430 418350
rect 21498 418294 21554 418350
rect 21622 418294 21678 418350
rect 21250 418170 21306 418226
rect 21374 418170 21430 418226
rect 21498 418170 21554 418226
rect 21622 418170 21678 418226
rect 21250 418046 21306 418102
rect 21374 418046 21430 418102
rect 21498 418046 21554 418102
rect 21622 418046 21678 418102
rect 21250 417922 21306 417978
rect 21374 417922 21430 417978
rect 21498 417922 21554 417978
rect 21622 417922 21678 417978
rect 21250 400294 21306 400350
rect 21374 400294 21430 400350
rect 21498 400294 21554 400350
rect 21622 400294 21678 400350
rect 21250 400170 21306 400226
rect 21374 400170 21430 400226
rect 21498 400170 21554 400226
rect 21622 400170 21678 400226
rect 21250 400046 21306 400102
rect 21374 400046 21430 400102
rect 21498 400046 21554 400102
rect 21622 400046 21678 400102
rect 21250 399922 21306 399978
rect 21374 399922 21430 399978
rect 21498 399922 21554 399978
rect 21622 399922 21678 399978
rect 21250 382294 21306 382350
rect 21374 382294 21430 382350
rect 21498 382294 21554 382350
rect 21622 382294 21678 382350
rect 21250 382170 21306 382226
rect 21374 382170 21430 382226
rect 21498 382170 21554 382226
rect 21622 382170 21678 382226
rect 21250 382046 21306 382102
rect 21374 382046 21430 382102
rect 21498 382046 21554 382102
rect 21622 382046 21678 382102
rect 21250 381922 21306 381978
rect 21374 381922 21430 381978
rect 21498 381922 21554 381978
rect 21622 381922 21678 381978
rect 21250 364294 21306 364350
rect 21374 364294 21430 364350
rect 21498 364294 21554 364350
rect 21622 364294 21678 364350
rect 21250 364170 21306 364226
rect 21374 364170 21430 364226
rect 21498 364170 21554 364226
rect 21622 364170 21678 364226
rect 21250 364046 21306 364102
rect 21374 364046 21430 364102
rect 21498 364046 21554 364102
rect 21622 364046 21678 364102
rect 21250 363922 21306 363978
rect 21374 363922 21430 363978
rect 21498 363922 21554 363978
rect 21622 363922 21678 363978
rect 21250 346294 21306 346350
rect 21374 346294 21430 346350
rect 21498 346294 21554 346350
rect 21622 346294 21678 346350
rect 21250 346170 21306 346226
rect 21374 346170 21430 346226
rect 21498 346170 21554 346226
rect 21622 346170 21678 346226
rect 21250 346046 21306 346102
rect 21374 346046 21430 346102
rect 21498 346046 21554 346102
rect 21622 346046 21678 346102
rect 21250 345922 21306 345978
rect 21374 345922 21430 345978
rect 21498 345922 21554 345978
rect 21622 345922 21678 345978
rect 21250 328294 21306 328350
rect 21374 328294 21430 328350
rect 21498 328294 21554 328350
rect 21622 328294 21678 328350
rect 21250 328170 21306 328226
rect 21374 328170 21430 328226
rect 21498 328170 21554 328226
rect 21622 328170 21678 328226
rect 21250 328046 21306 328102
rect 21374 328046 21430 328102
rect 21498 328046 21554 328102
rect 21622 328046 21678 328102
rect 21250 327922 21306 327978
rect 21374 327922 21430 327978
rect 21498 327922 21554 327978
rect 21622 327922 21678 327978
rect 21250 310294 21306 310350
rect 21374 310294 21430 310350
rect 21498 310294 21554 310350
rect 21622 310294 21678 310350
rect 21250 310170 21306 310226
rect 21374 310170 21430 310226
rect 21498 310170 21554 310226
rect 21622 310170 21678 310226
rect 21250 310046 21306 310102
rect 21374 310046 21430 310102
rect 21498 310046 21554 310102
rect 21622 310046 21678 310102
rect 21250 309922 21306 309978
rect 21374 309922 21430 309978
rect 21498 309922 21554 309978
rect 21622 309922 21678 309978
rect 21250 292294 21306 292350
rect 21374 292294 21430 292350
rect 21498 292294 21554 292350
rect 21622 292294 21678 292350
rect 21250 292170 21306 292226
rect 21374 292170 21430 292226
rect 21498 292170 21554 292226
rect 21622 292170 21678 292226
rect 21250 292046 21306 292102
rect 21374 292046 21430 292102
rect 21498 292046 21554 292102
rect 21622 292046 21678 292102
rect 21250 291922 21306 291978
rect 21374 291922 21430 291978
rect 21498 291922 21554 291978
rect 21622 291922 21678 291978
rect 21250 274294 21306 274350
rect 21374 274294 21430 274350
rect 21498 274294 21554 274350
rect 21622 274294 21678 274350
rect 21250 274170 21306 274226
rect 21374 274170 21430 274226
rect 21498 274170 21554 274226
rect 21622 274170 21678 274226
rect 21250 274046 21306 274102
rect 21374 274046 21430 274102
rect 21498 274046 21554 274102
rect 21622 274046 21678 274102
rect 21250 273922 21306 273978
rect 21374 273922 21430 273978
rect 21498 273922 21554 273978
rect 21622 273922 21678 273978
rect 21250 256294 21306 256350
rect 21374 256294 21430 256350
rect 21498 256294 21554 256350
rect 21622 256294 21678 256350
rect 21250 256170 21306 256226
rect 21374 256170 21430 256226
rect 21498 256170 21554 256226
rect 21622 256170 21678 256226
rect 21250 256046 21306 256102
rect 21374 256046 21430 256102
rect 21498 256046 21554 256102
rect 21622 256046 21678 256102
rect 21250 255922 21306 255978
rect 21374 255922 21430 255978
rect 21498 255922 21554 255978
rect 21622 255922 21678 255978
rect 21250 238294 21306 238350
rect 21374 238294 21430 238350
rect 21498 238294 21554 238350
rect 21622 238294 21678 238350
rect 21250 238170 21306 238226
rect 21374 238170 21430 238226
rect 21498 238170 21554 238226
rect 21622 238170 21678 238226
rect 21250 238046 21306 238102
rect 21374 238046 21430 238102
rect 21498 238046 21554 238102
rect 21622 238046 21678 238102
rect 21250 237922 21306 237978
rect 21374 237922 21430 237978
rect 21498 237922 21554 237978
rect 21622 237922 21678 237978
rect 21250 220294 21306 220350
rect 21374 220294 21430 220350
rect 21498 220294 21554 220350
rect 21622 220294 21678 220350
rect 21250 220170 21306 220226
rect 21374 220170 21430 220226
rect 21498 220170 21554 220226
rect 21622 220170 21678 220226
rect 21250 220046 21306 220102
rect 21374 220046 21430 220102
rect 21498 220046 21554 220102
rect 21622 220046 21678 220102
rect 21250 219922 21306 219978
rect 21374 219922 21430 219978
rect 21498 219922 21554 219978
rect 21622 219922 21678 219978
rect 21250 202294 21306 202350
rect 21374 202294 21430 202350
rect 21498 202294 21554 202350
rect 21622 202294 21678 202350
rect 21250 202170 21306 202226
rect 21374 202170 21430 202226
rect 21498 202170 21554 202226
rect 21622 202170 21678 202226
rect 21250 202046 21306 202102
rect 21374 202046 21430 202102
rect 21498 202046 21554 202102
rect 21622 202046 21678 202102
rect 21250 201922 21306 201978
rect 21374 201922 21430 201978
rect 21498 201922 21554 201978
rect 21622 201922 21678 201978
rect 21250 184294 21306 184350
rect 21374 184294 21430 184350
rect 21498 184294 21554 184350
rect 21622 184294 21678 184350
rect 21250 184170 21306 184226
rect 21374 184170 21430 184226
rect 21498 184170 21554 184226
rect 21622 184170 21678 184226
rect 21250 184046 21306 184102
rect 21374 184046 21430 184102
rect 21498 184046 21554 184102
rect 21622 184046 21678 184102
rect 21250 183922 21306 183978
rect 21374 183922 21430 183978
rect 21498 183922 21554 183978
rect 21622 183922 21678 183978
rect 21250 166294 21306 166350
rect 21374 166294 21430 166350
rect 21498 166294 21554 166350
rect 21622 166294 21678 166350
rect 21250 166170 21306 166226
rect 21374 166170 21430 166226
rect 21498 166170 21554 166226
rect 21622 166170 21678 166226
rect 21250 166046 21306 166102
rect 21374 166046 21430 166102
rect 21498 166046 21554 166102
rect 21622 166046 21678 166102
rect 21250 165922 21306 165978
rect 21374 165922 21430 165978
rect 21498 165922 21554 165978
rect 21622 165922 21678 165978
rect 21250 148294 21306 148350
rect 21374 148294 21430 148350
rect 21498 148294 21554 148350
rect 21622 148294 21678 148350
rect 21250 148170 21306 148226
rect 21374 148170 21430 148226
rect 21498 148170 21554 148226
rect 21622 148170 21678 148226
rect 21250 148046 21306 148102
rect 21374 148046 21430 148102
rect 21498 148046 21554 148102
rect 21622 148046 21678 148102
rect 21250 147922 21306 147978
rect 21374 147922 21430 147978
rect 21498 147922 21554 147978
rect 21622 147922 21678 147978
rect 21250 130294 21306 130350
rect 21374 130294 21430 130350
rect 21498 130294 21554 130350
rect 21622 130294 21678 130350
rect 21250 130170 21306 130226
rect 21374 130170 21430 130226
rect 21498 130170 21554 130226
rect 21622 130170 21678 130226
rect 21250 130046 21306 130102
rect 21374 130046 21430 130102
rect 21498 130046 21554 130102
rect 21622 130046 21678 130102
rect 21250 129922 21306 129978
rect 21374 129922 21430 129978
rect 21498 129922 21554 129978
rect 21622 129922 21678 129978
rect 21250 112294 21306 112350
rect 21374 112294 21430 112350
rect 21498 112294 21554 112350
rect 21622 112294 21678 112350
rect 21250 112170 21306 112226
rect 21374 112170 21430 112226
rect 21498 112170 21554 112226
rect 21622 112170 21678 112226
rect 21250 112046 21306 112102
rect 21374 112046 21430 112102
rect 21498 112046 21554 112102
rect 21622 112046 21678 112102
rect 21250 111922 21306 111978
rect 21374 111922 21430 111978
rect 21498 111922 21554 111978
rect 21622 111922 21678 111978
rect 21250 94294 21306 94350
rect 21374 94294 21430 94350
rect 21498 94294 21554 94350
rect 21622 94294 21678 94350
rect 21250 94170 21306 94226
rect 21374 94170 21430 94226
rect 21498 94170 21554 94226
rect 21622 94170 21678 94226
rect 21250 94046 21306 94102
rect 21374 94046 21430 94102
rect 21498 94046 21554 94102
rect 21622 94046 21678 94102
rect 21250 93922 21306 93978
rect 21374 93922 21430 93978
rect 21498 93922 21554 93978
rect 21622 93922 21678 93978
rect 21250 76294 21306 76350
rect 21374 76294 21430 76350
rect 21498 76294 21554 76350
rect 21622 76294 21678 76350
rect 21250 76170 21306 76226
rect 21374 76170 21430 76226
rect 21498 76170 21554 76226
rect 21622 76170 21678 76226
rect 21250 76046 21306 76102
rect 21374 76046 21430 76102
rect 21498 76046 21554 76102
rect 21622 76046 21678 76102
rect 21250 75922 21306 75978
rect 21374 75922 21430 75978
rect 21498 75922 21554 75978
rect 21622 75922 21678 75978
rect 21250 58294 21306 58350
rect 21374 58294 21430 58350
rect 21498 58294 21554 58350
rect 21622 58294 21678 58350
rect 21250 58170 21306 58226
rect 21374 58170 21430 58226
rect 21498 58170 21554 58226
rect 21622 58170 21678 58226
rect 21250 58046 21306 58102
rect 21374 58046 21430 58102
rect 21498 58046 21554 58102
rect 21622 58046 21678 58102
rect 21250 57922 21306 57978
rect 21374 57922 21430 57978
rect 21498 57922 21554 57978
rect 21622 57922 21678 57978
rect 21250 40294 21306 40350
rect 21374 40294 21430 40350
rect 21498 40294 21554 40350
rect 21622 40294 21678 40350
rect 21250 40170 21306 40226
rect 21374 40170 21430 40226
rect 21498 40170 21554 40226
rect 21622 40170 21678 40226
rect 21250 40046 21306 40102
rect 21374 40046 21430 40102
rect 21498 40046 21554 40102
rect 21622 40046 21678 40102
rect 21250 39922 21306 39978
rect 21374 39922 21430 39978
rect 21498 39922 21554 39978
rect 21622 39922 21678 39978
rect 21250 22294 21306 22350
rect 21374 22294 21430 22350
rect 21498 22294 21554 22350
rect 21622 22294 21678 22350
rect 21250 22170 21306 22226
rect 21374 22170 21430 22226
rect 21498 22170 21554 22226
rect 21622 22170 21678 22226
rect 21250 22046 21306 22102
rect 21374 22046 21430 22102
rect 21498 22046 21554 22102
rect 21622 22046 21678 22102
rect 21250 21922 21306 21978
rect 21374 21922 21430 21978
rect 21498 21922 21554 21978
rect 21622 21922 21678 21978
rect 21250 4294 21306 4350
rect 21374 4294 21430 4350
rect 21498 4294 21554 4350
rect 21622 4294 21678 4350
rect 21250 4170 21306 4226
rect 21374 4170 21430 4226
rect 21498 4170 21554 4226
rect 21622 4170 21678 4226
rect 21250 4046 21306 4102
rect 21374 4046 21430 4102
rect 21498 4046 21554 4102
rect 21622 4046 21678 4102
rect 21250 3922 21306 3978
rect 21374 3922 21430 3978
rect 21498 3922 21554 3978
rect 21622 3922 21678 3978
rect 21250 -216 21306 -160
rect 21374 -216 21430 -160
rect 21498 -216 21554 -160
rect 21622 -216 21678 -160
rect 21250 -340 21306 -284
rect 21374 -340 21430 -284
rect 21498 -340 21554 -284
rect 21622 -340 21678 -284
rect 21250 -464 21306 -408
rect 21374 -464 21430 -408
rect 21498 -464 21554 -408
rect 21622 -464 21678 -408
rect 21250 -588 21306 -532
rect 21374 -588 21430 -532
rect 21498 -588 21554 -532
rect 21622 -588 21678 -532
rect 24970 598116 25026 598172
rect 25094 598116 25150 598172
rect 25218 598116 25274 598172
rect 25342 598116 25398 598172
rect 24970 597992 25026 598048
rect 25094 597992 25150 598048
rect 25218 597992 25274 598048
rect 25342 597992 25398 598048
rect 24970 597868 25026 597924
rect 25094 597868 25150 597924
rect 25218 597868 25274 597924
rect 25342 597868 25398 597924
rect 24970 597744 25026 597800
rect 25094 597744 25150 597800
rect 25218 597744 25274 597800
rect 25342 597744 25398 597800
rect 24970 586294 25026 586350
rect 25094 586294 25150 586350
rect 25218 586294 25274 586350
rect 25342 586294 25398 586350
rect 24970 586170 25026 586226
rect 25094 586170 25150 586226
rect 25218 586170 25274 586226
rect 25342 586170 25398 586226
rect 24970 586046 25026 586102
rect 25094 586046 25150 586102
rect 25218 586046 25274 586102
rect 25342 586046 25398 586102
rect 24970 585922 25026 585978
rect 25094 585922 25150 585978
rect 25218 585922 25274 585978
rect 25342 585922 25398 585978
rect 24970 568294 25026 568350
rect 25094 568294 25150 568350
rect 25218 568294 25274 568350
rect 25342 568294 25398 568350
rect 24970 568170 25026 568226
rect 25094 568170 25150 568226
rect 25218 568170 25274 568226
rect 25342 568170 25398 568226
rect 24970 568046 25026 568102
rect 25094 568046 25150 568102
rect 25218 568046 25274 568102
rect 25342 568046 25398 568102
rect 24970 567922 25026 567978
rect 25094 567922 25150 567978
rect 25218 567922 25274 567978
rect 25342 567922 25398 567978
rect 24970 550294 25026 550350
rect 25094 550294 25150 550350
rect 25218 550294 25274 550350
rect 25342 550294 25398 550350
rect 24970 550170 25026 550226
rect 25094 550170 25150 550226
rect 25218 550170 25274 550226
rect 25342 550170 25398 550226
rect 24970 550046 25026 550102
rect 25094 550046 25150 550102
rect 25218 550046 25274 550102
rect 25342 550046 25398 550102
rect 24970 549922 25026 549978
rect 25094 549922 25150 549978
rect 25218 549922 25274 549978
rect 25342 549922 25398 549978
rect 24970 532294 25026 532350
rect 25094 532294 25150 532350
rect 25218 532294 25274 532350
rect 25342 532294 25398 532350
rect 24970 532170 25026 532226
rect 25094 532170 25150 532226
rect 25218 532170 25274 532226
rect 25342 532170 25398 532226
rect 24970 532046 25026 532102
rect 25094 532046 25150 532102
rect 25218 532046 25274 532102
rect 25342 532046 25398 532102
rect 24970 531922 25026 531978
rect 25094 531922 25150 531978
rect 25218 531922 25274 531978
rect 25342 531922 25398 531978
rect 24970 514294 25026 514350
rect 25094 514294 25150 514350
rect 25218 514294 25274 514350
rect 25342 514294 25398 514350
rect 24970 514170 25026 514226
rect 25094 514170 25150 514226
rect 25218 514170 25274 514226
rect 25342 514170 25398 514226
rect 24970 514046 25026 514102
rect 25094 514046 25150 514102
rect 25218 514046 25274 514102
rect 25342 514046 25398 514102
rect 24970 513922 25026 513978
rect 25094 513922 25150 513978
rect 25218 513922 25274 513978
rect 25342 513922 25398 513978
rect 24970 496294 25026 496350
rect 25094 496294 25150 496350
rect 25218 496294 25274 496350
rect 25342 496294 25398 496350
rect 24970 496170 25026 496226
rect 25094 496170 25150 496226
rect 25218 496170 25274 496226
rect 25342 496170 25398 496226
rect 24970 496046 25026 496102
rect 25094 496046 25150 496102
rect 25218 496046 25274 496102
rect 25342 496046 25398 496102
rect 24970 495922 25026 495978
rect 25094 495922 25150 495978
rect 25218 495922 25274 495978
rect 25342 495922 25398 495978
rect 24970 478294 25026 478350
rect 25094 478294 25150 478350
rect 25218 478294 25274 478350
rect 25342 478294 25398 478350
rect 24970 478170 25026 478226
rect 25094 478170 25150 478226
rect 25218 478170 25274 478226
rect 25342 478170 25398 478226
rect 24970 478046 25026 478102
rect 25094 478046 25150 478102
rect 25218 478046 25274 478102
rect 25342 478046 25398 478102
rect 24970 477922 25026 477978
rect 25094 477922 25150 477978
rect 25218 477922 25274 477978
rect 25342 477922 25398 477978
rect 24970 460294 25026 460350
rect 25094 460294 25150 460350
rect 25218 460294 25274 460350
rect 25342 460294 25398 460350
rect 24970 460170 25026 460226
rect 25094 460170 25150 460226
rect 25218 460170 25274 460226
rect 25342 460170 25398 460226
rect 24970 460046 25026 460102
rect 25094 460046 25150 460102
rect 25218 460046 25274 460102
rect 25342 460046 25398 460102
rect 24970 459922 25026 459978
rect 25094 459922 25150 459978
rect 25218 459922 25274 459978
rect 25342 459922 25398 459978
rect 24970 442294 25026 442350
rect 25094 442294 25150 442350
rect 25218 442294 25274 442350
rect 25342 442294 25398 442350
rect 24970 442170 25026 442226
rect 25094 442170 25150 442226
rect 25218 442170 25274 442226
rect 25342 442170 25398 442226
rect 24970 442046 25026 442102
rect 25094 442046 25150 442102
rect 25218 442046 25274 442102
rect 25342 442046 25398 442102
rect 24970 441922 25026 441978
rect 25094 441922 25150 441978
rect 25218 441922 25274 441978
rect 25342 441922 25398 441978
rect 24970 424294 25026 424350
rect 25094 424294 25150 424350
rect 25218 424294 25274 424350
rect 25342 424294 25398 424350
rect 24970 424170 25026 424226
rect 25094 424170 25150 424226
rect 25218 424170 25274 424226
rect 25342 424170 25398 424226
rect 24970 424046 25026 424102
rect 25094 424046 25150 424102
rect 25218 424046 25274 424102
rect 25342 424046 25398 424102
rect 24970 423922 25026 423978
rect 25094 423922 25150 423978
rect 25218 423922 25274 423978
rect 25342 423922 25398 423978
rect 24970 406294 25026 406350
rect 25094 406294 25150 406350
rect 25218 406294 25274 406350
rect 25342 406294 25398 406350
rect 24970 406170 25026 406226
rect 25094 406170 25150 406226
rect 25218 406170 25274 406226
rect 25342 406170 25398 406226
rect 24970 406046 25026 406102
rect 25094 406046 25150 406102
rect 25218 406046 25274 406102
rect 25342 406046 25398 406102
rect 24970 405922 25026 405978
rect 25094 405922 25150 405978
rect 25218 405922 25274 405978
rect 25342 405922 25398 405978
rect 24970 388294 25026 388350
rect 25094 388294 25150 388350
rect 25218 388294 25274 388350
rect 25342 388294 25398 388350
rect 24970 388170 25026 388226
rect 25094 388170 25150 388226
rect 25218 388170 25274 388226
rect 25342 388170 25398 388226
rect 24970 388046 25026 388102
rect 25094 388046 25150 388102
rect 25218 388046 25274 388102
rect 25342 388046 25398 388102
rect 24970 387922 25026 387978
rect 25094 387922 25150 387978
rect 25218 387922 25274 387978
rect 25342 387922 25398 387978
rect 24970 370294 25026 370350
rect 25094 370294 25150 370350
rect 25218 370294 25274 370350
rect 25342 370294 25398 370350
rect 24970 370170 25026 370226
rect 25094 370170 25150 370226
rect 25218 370170 25274 370226
rect 25342 370170 25398 370226
rect 24970 370046 25026 370102
rect 25094 370046 25150 370102
rect 25218 370046 25274 370102
rect 25342 370046 25398 370102
rect 24970 369922 25026 369978
rect 25094 369922 25150 369978
rect 25218 369922 25274 369978
rect 25342 369922 25398 369978
rect 24970 352294 25026 352350
rect 25094 352294 25150 352350
rect 25218 352294 25274 352350
rect 25342 352294 25398 352350
rect 24970 352170 25026 352226
rect 25094 352170 25150 352226
rect 25218 352170 25274 352226
rect 25342 352170 25398 352226
rect 24970 352046 25026 352102
rect 25094 352046 25150 352102
rect 25218 352046 25274 352102
rect 25342 352046 25398 352102
rect 24970 351922 25026 351978
rect 25094 351922 25150 351978
rect 25218 351922 25274 351978
rect 25342 351922 25398 351978
rect 24970 334294 25026 334350
rect 25094 334294 25150 334350
rect 25218 334294 25274 334350
rect 25342 334294 25398 334350
rect 24970 334170 25026 334226
rect 25094 334170 25150 334226
rect 25218 334170 25274 334226
rect 25342 334170 25398 334226
rect 24970 334046 25026 334102
rect 25094 334046 25150 334102
rect 25218 334046 25274 334102
rect 25342 334046 25398 334102
rect 24970 333922 25026 333978
rect 25094 333922 25150 333978
rect 25218 333922 25274 333978
rect 25342 333922 25398 333978
rect 24970 316294 25026 316350
rect 25094 316294 25150 316350
rect 25218 316294 25274 316350
rect 25342 316294 25398 316350
rect 24970 316170 25026 316226
rect 25094 316170 25150 316226
rect 25218 316170 25274 316226
rect 25342 316170 25398 316226
rect 24970 316046 25026 316102
rect 25094 316046 25150 316102
rect 25218 316046 25274 316102
rect 25342 316046 25398 316102
rect 24970 315922 25026 315978
rect 25094 315922 25150 315978
rect 25218 315922 25274 315978
rect 25342 315922 25398 315978
rect 24970 298294 25026 298350
rect 25094 298294 25150 298350
rect 25218 298294 25274 298350
rect 25342 298294 25398 298350
rect 24970 298170 25026 298226
rect 25094 298170 25150 298226
rect 25218 298170 25274 298226
rect 25342 298170 25398 298226
rect 24970 298046 25026 298102
rect 25094 298046 25150 298102
rect 25218 298046 25274 298102
rect 25342 298046 25398 298102
rect 24970 297922 25026 297978
rect 25094 297922 25150 297978
rect 25218 297922 25274 297978
rect 25342 297922 25398 297978
rect 24970 280294 25026 280350
rect 25094 280294 25150 280350
rect 25218 280294 25274 280350
rect 25342 280294 25398 280350
rect 24970 280170 25026 280226
rect 25094 280170 25150 280226
rect 25218 280170 25274 280226
rect 25342 280170 25398 280226
rect 24970 280046 25026 280102
rect 25094 280046 25150 280102
rect 25218 280046 25274 280102
rect 25342 280046 25398 280102
rect 24970 279922 25026 279978
rect 25094 279922 25150 279978
rect 25218 279922 25274 279978
rect 25342 279922 25398 279978
rect 24970 262294 25026 262350
rect 25094 262294 25150 262350
rect 25218 262294 25274 262350
rect 25342 262294 25398 262350
rect 24970 262170 25026 262226
rect 25094 262170 25150 262226
rect 25218 262170 25274 262226
rect 25342 262170 25398 262226
rect 24970 262046 25026 262102
rect 25094 262046 25150 262102
rect 25218 262046 25274 262102
rect 25342 262046 25398 262102
rect 24970 261922 25026 261978
rect 25094 261922 25150 261978
rect 25218 261922 25274 261978
rect 25342 261922 25398 261978
rect 24970 244294 25026 244350
rect 25094 244294 25150 244350
rect 25218 244294 25274 244350
rect 25342 244294 25398 244350
rect 24970 244170 25026 244226
rect 25094 244170 25150 244226
rect 25218 244170 25274 244226
rect 25342 244170 25398 244226
rect 24970 244046 25026 244102
rect 25094 244046 25150 244102
rect 25218 244046 25274 244102
rect 25342 244046 25398 244102
rect 24970 243922 25026 243978
rect 25094 243922 25150 243978
rect 25218 243922 25274 243978
rect 25342 243922 25398 243978
rect 24970 226294 25026 226350
rect 25094 226294 25150 226350
rect 25218 226294 25274 226350
rect 25342 226294 25398 226350
rect 24970 226170 25026 226226
rect 25094 226170 25150 226226
rect 25218 226170 25274 226226
rect 25342 226170 25398 226226
rect 24970 226046 25026 226102
rect 25094 226046 25150 226102
rect 25218 226046 25274 226102
rect 25342 226046 25398 226102
rect 24970 225922 25026 225978
rect 25094 225922 25150 225978
rect 25218 225922 25274 225978
rect 25342 225922 25398 225978
rect 24970 208294 25026 208350
rect 25094 208294 25150 208350
rect 25218 208294 25274 208350
rect 25342 208294 25398 208350
rect 24970 208170 25026 208226
rect 25094 208170 25150 208226
rect 25218 208170 25274 208226
rect 25342 208170 25398 208226
rect 24970 208046 25026 208102
rect 25094 208046 25150 208102
rect 25218 208046 25274 208102
rect 25342 208046 25398 208102
rect 24970 207922 25026 207978
rect 25094 207922 25150 207978
rect 25218 207922 25274 207978
rect 25342 207922 25398 207978
rect 24970 190294 25026 190350
rect 25094 190294 25150 190350
rect 25218 190294 25274 190350
rect 25342 190294 25398 190350
rect 24970 190170 25026 190226
rect 25094 190170 25150 190226
rect 25218 190170 25274 190226
rect 25342 190170 25398 190226
rect 24970 190046 25026 190102
rect 25094 190046 25150 190102
rect 25218 190046 25274 190102
rect 25342 190046 25398 190102
rect 24970 189922 25026 189978
rect 25094 189922 25150 189978
rect 25218 189922 25274 189978
rect 25342 189922 25398 189978
rect 24970 172294 25026 172350
rect 25094 172294 25150 172350
rect 25218 172294 25274 172350
rect 25342 172294 25398 172350
rect 24970 172170 25026 172226
rect 25094 172170 25150 172226
rect 25218 172170 25274 172226
rect 25342 172170 25398 172226
rect 24970 172046 25026 172102
rect 25094 172046 25150 172102
rect 25218 172046 25274 172102
rect 25342 172046 25398 172102
rect 24970 171922 25026 171978
rect 25094 171922 25150 171978
rect 25218 171922 25274 171978
rect 25342 171922 25398 171978
rect 24970 154294 25026 154350
rect 25094 154294 25150 154350
rect 25218 154294 25274 154350
rect 25342 154294 25398 154350
rect 24970 154170 25026 154226
rect 25094 154170 25150 154226
rect 25218 154170 25274 154226
rect 25342 154170 25398 154226
rect 24970 154046 25026 154102
rect 25094 154046 25150 154102
rect 25218 154046 25274 154102
rect 25342 154046 25398 154102
rect 24970 153922 25026 153978
rect 25094 153922 25150 153978
rect 25218 153922 25274 153978
rect 25342 153922 25398 153978
rect 24970 136294 25026 136350
rect 25094 136294 25150 136350
rect 25218 136294 25274 136350
rect 25342 136294 25398 136350
rect 24970 136170 25026 136226
rect 25094 136170 25150 136226
rect 25218 136170 25274 136226
rect 25342 136170 25398 136226
rect 24970 136046 25026 136102
rect 25094 136046 25150 136102
rect 25218 136046 25274 136102
rect 25342 136046 25398 136102
rect 24970 135922 25026 135978
rect 25094 135922 25150 135978
rect 25218 135922 25274 135978
rect 25342 135922 25398 135978
rect 24970 118294 25026 118350
rect 25094 118294 25150 118350
rect 25218 118294 25274 118350
rect 25342 118294 25398 118350
rect 24970 118170 25026 118226
rect 25094 118170 25150 118226
rect 25218 118170 25274 118226
rect 25342 118170 25398 118226
rect 24970 118046 25026 118102
rect 25094 118046 25150 118102
rect 25218 118046 25274 118102
rect 25342 118046 25398 118102
rect 24970 117922 25026 117978
rect 25094 117922 25150 117978
rect 25218 117922 25274 117978
rect 25342 117922 25398 117978
rect 24970 100294 25026 100350
rect 25094 100294 25150 100350
rect 25218 100294 25274 100350
rect 25342 100294 25398 100350
rect 24970 100170 25026 100226
rect 25094 100170 25150 100226
rect 25218 100170 25274 100226
rect 25342 100170 25398 100226
rect 24970 100046 25026 100102
rect 25094 100046 25150 100102
rect 25218 100046 25274 100102
rect 25342 100046 25398 100102
rect 24970 99922 25026 99978
rect 25094 99922 25150 99978
rect 25218 99922 25274 99978
rect 25342 99922 25398 99978
rect 24970 82294 25026 82350
rect 25094 82294 25150 82350
rect 25218 82294 25274 82350
rect 25342 82294 25398 82350
rect 24970 82170 25026 82226
rect 25094 82170 25150 82226
rect 25218 82170 25274 82226
rect 25342 82170 25398 82226
rect 24970 82046 25026 82102
rect 25094 82046 25150 82102
rect 25218 82046 25274 82102
rect 25342 82046 25398 82102
rect 24970 81922 25026 81978
rect 25094 81922 25150 81978
rect 25218 81922 25274 81978
rect 25342 81922 25398 81978
rect 24970 64294 25026 64350
rect 25094 64294 25150 64350
rect 25218 64294 25274 64350
rect 25342 64294 25398 64350
rect 24970 64170 25026 64226
rect 25094 64170 25150 64226
rect 25218 64170 25274 64226
rect 25342 64170 25398 64226
rect 24970 64046 25026 64102
rect 25094 64046 25150 64102
rect 25218 64046 25274 64102
rect 25342 64046 25398 64102
rect 24970 63922 25026 63978
rect 25094 63922 25150 63978
rect 25218 63922 25274 63978
rect 25342 63922 25398 63978
rect 24970 46294 25026 46350
rect 25094 46294 25150 46350
rect 25218 46294 25274 46350
rect 25342 46294 25398 46350
rect 24970 46170 25026 46226
rect 25094 46170 25150 46226
rect 25218 46170 25274 46226
rect 25342 46170 25398 46226
rect 24970 46046 25026 46102
rect 25094 46046 25150 46102
rect 25218 46046 25274 46102
rect 25342 46046 25398 46102
rect 24970 45922 25026 45978
rect 25094 45922 25150 45978
rect 25218 45922 25274 45978
rect 25342 45922 25398 45978
rect 24970 28294 25026 28350
rect 25094 28294 25150 28350
rect 25218 28294 25274 28350
rect 25342 28294 25398 28350
rect 24970 28170 25026 28226
rect 25094 28170 25150 28226
rect 25218 28170 25274 28226
rect 25342 28170 25398 28226
rect 24970 28046 25026 28102
rect 25094 28046 25150 28102
rect 25218 28046 25274 28102
rect 25342 28046 25398 28102
rect 24970 27922 25026 27978
rect 25094 27922 25150 27978
rect 25218 27922 25274 27978
rect 25342 27922 25398 27978
rect 24970 10294 25026 10350
rect 25094 10294 25150 10350
rect 25218 10294 25274 10350
rect 25342 10294 25398 10350
rect 24970 10170 25026 10226
rect 25094 10170 25150 10226
rect 25218 10170 25274 10226
rect 25342 10170 25398 10226
rect 24970 10046 25026 10102
rect 25094 10046 25150 10102
rect 25218 10046 25274 10102
rect 25342 10046 25398 10102
rect 24970 9922 25026 9978
rect 25094 9922 25150 9978
rect 25218 9922 25274 9978
rect 25342 9922 25398 9978
rect 24970 -1176 25026 -1120
rect 25094 -1176 25150 -1120
rect 25218 -1176 25274 -1120
rect 25342 -1176 25398 -1120
rect 24970 -1300 25026 -1244
rect 25094 -1300 25150 -1244
rect 25218 -1300 25274 -1244
rect 25342 -1300 25398 -1244
rect 24970 -1424 25026 -1368
rect 25094 -1424 25150 -1368
rect 25218 -1424 25274 -1368
rect 25342 -1424 25398 -1368
rect 24970 -1548 25026 -1492
rect 25094 -1548 25150 -1492
rect 25218 -1548 25274 -1492
rect 25342 -1548 25398 -1492
rect 39250 597156 39306 597212
rect 39374 597156 39430 597212
rect 39498 597156 39554 597212
rect 39622 597156 39678 597212
rect 39250 597032 39306 597088
rect 39374 597032 39430 597088
rect 39498 597032 39554 597088
rect 39622 597032 39678 597088
rect 39250 596908 39306 596964
rect 39374 596908 39430 596964
rect 39498 596908 39554 596964
rect 39622 596908 39678 596964
rect 39250 596784 39306 596840
rect 39374 596784 39430 596840
rect 39498 596784 39554 596840
rect 39622 596784 39678 596840
rect 39250 580294 39306 580350
rect 39374 580294 39430 580350
rect 39498 580294 39554 580350
rect 39622 580294 39678 580350
rect 39250 580170 39306 580226
rect 39374 580170 39430 580226
rect 39498 580170 39554 580226
rect 39622 580170 39678 580226
rect 39250 580046 39306 580102
rect 39374 580046 39430 580102
rect 39498 580046 39554 580102
rect 39622 580046 39678 580102
rect 39250 579922 39306 579978
rect 39374 579922 39430 579978
rect 39498 579922 39554 579978
rect 39622 579922 39678 579978
rect 39250 562294 39306 562350
rect 39374 562294 39430 562350
rect 39498 562294 39554 562350
rect 39622 562294 39678 562350
rect 39250 562170 39306 562226
rect 39374 562170 39430 562226
rect 39498 562170 39554 562226
rect 39622 562170 39678 562226
rect 39250 562046 39306 562102
rect 39374 562046 39430 562102
rect 39498 562046 39554 562102
rect 39622 562046 39678 562102
rect 39250 561922 39306 561978
rect 39374 561922 39430 561978
rect 39498 561922 39554 561978
rect 39622 561922 39678 561978
rect 39250 544294 39306 544350
rect 39374 544294 39430 544350
rect 39498 544294 39554 544350
rect 39622 544294 39678 544350
rect 39250 544170 39306 544226
rect 39374 544170 39430 544226
rect 39498 544170 39554 544226
rect 39622 544170 39678 544226
rect 39250 544046 39306 544102
rect 39374 544046 39430 544102
rect 39498 544046 39554 544102
rect 39622 544046 39678 544102
rect 39250 543922 39306 543978
rect 39374 543922 39430 543978
rect 39498 543922 39554 543978
rect 39622 543922 39678 543978
rect 39250 526294 39306 526350
rect 39374 526294 39430 526350
rect 39498 526294 39554 526350
rect 39622 526294 39678 526350
rect 39250 526170 39306 526226
rect 39374 526170 39430 526226
rect 39498 526170 39554 526226
rect 39622 526170 39678 526226
rect 39250 526046 39306 526102
rect 39374 526046 39430 526102
rect 39498 526046 39554 526102
rect 39622 526046 39678 526102
rect 39250 525922 39306 525978
rect 39374 525922 39430 525978
rect 39498 525922 39554 525978
rect 39622 525922 39678 525978
rect 39250 508294 39306 508350
rect 39374 508294 39430 508350
rect 39498 508294 39554 508350
rect 39622 508294 39678 508350
rect 39250 508170 39306 508226
rect 39374 508170 39430 508226
rect 39498 508170 39554 508226
rect 39622 508170 39678 508226
rect 39250 508046 39306 508102
rect 39374 508046 39430 508102
rect 39498 508046 39554 508102
rect 39622 508046 39678 508102
rect 39250 507922 39306 507978
rect 39374 507922 39430 507978
rect 39498 507922 39554 507978
rect 39622 507922 39678 507978
rect 39250 490294 39306 490350
rect 39374 490294 39430 490350
rect 39498 490294 39554 490350
rect 39622 490294 39678 490350
rect 39250 490170 39306 490226
rect 39374 490170 39430 490226
rect 39498 490170 39554 490226
rect 39622 490170 39678 490226
rect 39250 490046 39306 490102
rect 39374 490046 39430 490102
rect 39498 490046 39554 490102
rect 39622 490046 39678 490102
rect 39250 489922 39306 489978
rect 39374 489922 39430 489978
rect 39498 489922 39554 489978
rect 39622 489922 39678 489978
rect 39250 472294 39306 472350
rect 39374 472294 39430 472350
rect 39498 472294 39554 472350
rect 39622 472294 39678 472350
rect 39250 472170 39306 472226
rect 39374 472170 39430 472226
rect 39498 472170 39554 472226
rect 39622 472170 39678 472226
rect 39250 472046 39306 472102
rect 39374 472046 39430 472102
rect 39498 472046 39554 472102
rect 39622 472046 39678 472102
rect 39250 471922 39306 471978
rect 39374 471922 39430 471978
rect 39498 471922 39554 471978
rect 39622 471922 39678 471978
rect 39250 454294 39306 454350
rect 39374 454294 39430 454350
rect 39498 454294 39554 454350
rect 39622 454294 39678 454350
rect 39250 454170 39306 454226
rect 39374 454170 39430 454226
rect 39498 454170 39554 454226
rect 39622 454170 39678 454226
rect 39250 454046 39306 454102
rect 39374 454046 39430 454102
rect 39498 454046 39554 454102
rect 39622 454046 39678 454102
rect 39250 453922 39306 453978
rect 39374 453922 39430 453978
rect 39498 453922 39554 453978
rect 39622 453922 39678 453978
rect 39250 436294 39306 436350
rect 39374 436294 39430 436350
rect 39498 436294 39554 436350
rect 39622 436294 39678 436350
rect 39250 436170 39306 436226
rect 39374 436170 39430 436226
rect 39498 436170 39554 436226
rect 39622 436170 39678 436226
rect 39250 436046 39306 436102
rect 39374 436046 39430 436102
rect 39498 436046 39554 436102
rect 39622 436046 39678 436102
rect 39250 435922 39306 435978
rect 39374 435922 39430 435978
rect 39498 435922 39554 435978
rect 39622 435922 39678 435978
rect 39250 418294 39306 418350
rect 39374 418294 39430 418350
rect 39498 418294 39554 418350
rect 39622 418294 39678 418350
rect 39250 418170 39306 418226
rect 39374 418170 39430 418226
rect 39498 418170 39554 418226
rect 39622 418170 39678 418226
rect 39250 418046 39306 418102
rect 39374 418046 39430 418102
rect 39498 418046 39554 418102
rect 39622 418046 39678 418102
rect 39250 417922 39306 417978
rect 39374 417922 39430 417978
rect 39498 417922 39554 417978
rect 39622 417922 39678 417978
rect 39250 400294 39306 400350
rect 39374 400294 39430 400350
rect 39498 400294 39554 400350
rect 39622 400294 39678 400350
rect 39250 400170 39306 400226
rect 39374 400170 39430 400226
rect 39498 400170 39554 400226
rect 39622 400170 39678 400226
rect 39250 400046 39306 400102
rect 39374 400046 39430 400102
rect 39498 400046 39554 400102
rect 39622 400046 39678 400102
rect 39250 399922 39306 399978
rect 39374 399922 39430 399978
rect 39498 399922 39554 399978
rect 39622 399922 39678 399978
rect 39250 382294 39306 382350
rect 39374 382294 39430 382350
rect 39498 382294 39554 382350
rect 39622 382294 39678 382350
rect 39250 382170 39306 382226
rect 39374 382170 39430 382226
rect 39498 382170 39554 382226
rect 39622 382170 39678 382226
rect 39250 382046 39306 382102
rect 39374 382046 39430 382102
rect 39498 382046 39554 382102
rect 39622 382046 39678 382102
rect 39250 381922 39306 381978
rect 39374 381922 39430 381978
rect 39498 381922 39554 381978
rect 39622 381922 39678 381978
rect 39250 364294 39306 364350
rect 39374 364294 39430 364350
rect 39498 364294 39554 364350
rect 39622 364294 39678 364350
rect 39250 364170 39306 364226
rect 39374 364170 39430 364226
rect 39498 364170 39554 364226
rect 39622 364170 39678 364226
rect 39250 364046 39306 364102
rect 39374 364046 39430 364102
rect 39498 364046 39554 364102
rect 39622 364046 39678 364102
rect 39250 363922 39306 363978
rect 39374 363922 39430 363978
rect 39498 363922 39554 363978
rect 39622 363922 39678 363978
rect 39250 346294 39306 346350
rect 39374 346294 39430 346350
rect 39498 346294 39554 346350
rect 39622 346294 39678 346350
rect 39250 346170 39306 346226
rect 39374 346170 39430 346226
rect 39498 346170 39554 346226
rect 39622 346170 39678 346226
rect 39250 346046 39306 346102
rect 39374 346046 39430 346102
rect 39498 346046 39554 346102
rect 39622 346046 39678 346102
rect 39250 345922 39306 345978
rect 39374 345922 39430 345978
rect 39498 345922 39554 345978
rect 39622 345922 39678 345978
rect 39250 328294 39306 328350
rect 39374 328294 39430 328350
rect 39498 328294 39554 328350
rect 39622 328294 39678 328350
rect 39250 328170 39306 328226
rect 39374 328170 39430 328226
rect 39498 328170 39554 328226
rect 39622 328170 39678 328226
rect 39250 328046 39306 328102
rect 39374 328046 39430 328102
rect 39498 328046 39554 328102
rect 39622 328046 39678 328102
rect 39250 327922 39306 327978
rect 39374 327922 39430 327978
rect 39498 327922 39554 327978
rect 39622 327922 39678 327978
rect 39250 310294 39306 310350
rect 39374 310294 39430 310350
rect 39498 310294 39554 310350
rect 39622 310294 39678 310350
rect 39250 310170 39306 310226
rect 39374 310170 39430 310226
rect 39498 310170 39554 310226
rect 39622 310170 39678 310226
rect 39250 310046 39306 310102
rect 39374 310046 39430 310102
rect 39498 310046 39554 310102
rect 39622 310046 39678 310102
rect 39250 309922 39306 309978
rect 39374 309922 39430 309978
rect 39498 309922 39554 309978
rect 39622 309922 39678 309978
rect 39250 292294 39306 292350
rect 39374 292294 39430 292350
rect 39498 292294 39554 292350
rect 39622 292294 39678 292350
rect 39250 292170 39306 292226
rect 39374 292170 39430 292226
rect 39498 292170 39554 292226
rect 39622 292170 39678 292226
rect 39250 292046 39306 292102
rect 39374 292046 39430 292102
rect 39498 292046 39554 292102
rect 39622 292046 39678 292102
rect 39250 291922 39306 291978
rect 39374 291922 39430 291978
rect 39498 291922 39554 291978
rect 39622 291922 39678 291978
rect 39250 274294 39306 274350
rect 39374 274294 39430 274350
rect 39498 274294 39554 274350
rect 39622 274294 39678 274350
rect 39250 274170 39306 274226
rect 39374 274170 39430 274226
rect 39498 274170 39554 274226
rect 39622 274170 39678 274226
rect 39250 274046 39306 274102
rect 39374 274046 39430 274102
rect 39498 274046 39554 274102
rect 39622 274046 39678 274102
rect 39250 273922 39306 273978
rect 39374 273922 39430 273978
rect 39498 273922 39554 273978
rect 39622 273922 39678 273978
rect 39250 256294 39306 256350
rect 39374 256294 39430 256350
rect 39498 256294 39554 256350
rect 39622 256294 39678 256350
rect 39250 256170 39306 256226
rect 39374 256170 39430 256226
rect 39498 256170 39554 256226
rect 39622 256170 39678 256226
rect 39250 256046 39306 256102
rect 39374 256046 39430 256102
rect 39498 256046 39554 256102
rect 39622 256046 39678 256102
rect 39250 255922 39306 255978
rect 39374 255922 39430 255978
rect 39498 255922 39554 255978
rect 39622 255922 39678 255978
rect 39250 238294 39306 238350
rect 39374 238294 39430 238350
rect 39498 238294 39554 238350
rect 39622 238294 39678 238350
rect 39250 238170 39306 238226
rect 39374 238170 39430 238226
rect 39498 238170 39554 238226
rect 39622 238170 39678 238226
rect 39250 238046 39306 238102
rect 39374 238046 39430 238102
rect 39498 238046 39554 238102
rect 39622 238046 39678 238102
rect 39250 237922 39306 237978
rect 39374 237922 39430 237978
rect 39498 237922 39554 237978
rect 39622 237922 39678 237978
rect 39250 220294 39306 220350
rect 39374 220294 39430 220350
rect 39498 220294 39554 220350
rect 39622 220294 39678 220350
rect 39250 220170 39306 220226
rect 39374 220170 39430 220226
rect 39498 220170 39554 220226
rect 39622 220170 39678 220226
rect 39250 220046 39306 220102
rect 39374 220046 39430 220102
rect 39498 220046 39554 220102
rect 39622 220046 39678 220102
rect 39250 219922 39306 219978
rect 39374 219922 39430 219978
rect 39498 219922 39554 219978
rect 39622 219922 39678 219978
rect 39250 202294 39306 202350
rect 39374 202294 39430 202350
rect 39498 202294 39554 202350
rect 39622 202294 39678 202350
rect 39250 202170 39306 202226
rect 39374 202170 39430 202226
rect 39498 202170 39554 202226
rect 39622 202170 39678 202226
rect 39250 202046 39306 202102
rect 39374 202046 39430 202102
rect 39498 202046 39554 202102
rect 39622 202046 39678 202102
rect 39250 201922 39306 201978
rect 39374 201922 39430 201978
rect 39498 201922 39554 201978
rect 39622 201922 39678 201978
rect 39250 184294 39306 184350
rect 39374 184294 39430 184350
rect 39498 184294 39554 184350
rect 39622 184294 39678 184350
rect 39250 184170 39306 184226
rect 39374 184170 39430 184226
rect 39498 184170 39554 184226
rect 39622 184170 39678 184226
rect 39250 184046 39306 184102
rect 39374 184046 39430 184102
rect 39498 184046 39554 184102
rect 39622 184046 39678 184102
rect 39250 183922 39306 183978
rect 39374 183922 39430 183978
rect 39498 183922 39554 183978
rect 39622 183922 39678 183978
rect 39250 166294 39306 166350
rect 39374 166294 39430 166350
rect 39498 166294 39554 166350
rect 39622 166294 39678 166350
rect 39250 166170 39306 166226
rect 39374 166170 39430 166226
rect 39498 166170 39554 166226
rect 39622 166170 39678 166226
rect 39250 166046 39306 166102
rect 39374 166046 39430 166102
rect 39498 166046 39554 166102
rect 39622 166046 39678 166102
rect 39250 165922 39306 165978
rect 39374 165922 39430 165978
rect 39498 165922 39554 165978
rect 39622 165922 39678 165978
rect 39250 148294 39306 148350
rect 39374 148294 39430 148350
rect 39498 148294 39554 148350
rect 39622 148294 39678 148350
rect 39250 148170 39306 148226
rect 39374 148170 39430 148226
rect 39498 148170 39554 148226
rect 39622 148170 39678 148226
rect 39250 148046 39306 148102
rect 39374 148046 39430 148102
rect 39498 148046 39554 148102
rect 39622 148046 39678 148102
rect 39250 147922 39306 147978
rect 39374 147922 39430 147978
rect 39498 147922 39554 147978
rect 39622 147922 39678 147978
rect 39250 130294 39306 130350
rect 39374 130294 39430 130350
rect 39498 130294 39554 130350
rect 39622 130294 39678 130350
rect 39250 130170 39306 130226
rect 39374 130170 39430 130226
rect 39498 130170 39554 130226
rect 39622 130170 39678 130226
rect 39250 130046 39306 130102
rect 39374 130046 39430 130102
rect 39498 130046 39554 130102
rect 39622 130046 39678 130102
rect 39250 129922 39306 129978
rect 39374 129922 39430 129978
rect 39498 129922 39554 129978
rect 39622 129922 39678 129978
rect 39250 112294 39306 112350
rect 39374 112294 39430 112350
rect 39498 112294 39554 112350
rect 39622 112294 39678 112350
rect 39250 112170 39306 112226
rect 39374 112170 39430 112226
rect 39498 112170 39554 112226
rect 39622 112170 39678 112226
rect 39250 112046 39306 112102
rect 39374 112046 39430 112102
rect 39498 112046 39554 112102
rect 39622 112046 39678 112102
rect 39250 111922 39306 111978
rect 39374 111922 39430 111978
rect 39498 111922 39554 111978
rect 39622 111922 39678 111978
rect 39250 94294 39306 94350
rect 39374 94294 39430 94350
rect 39498 94294 39554 94350
rect 39622 94294 39678 94350
rect 39250 94170 39306 94226
rect 39374 94170 39430 94226
rect 39498 94170 39554 94226
rect 39622 94170 39678 94226
rect 39250 94046 39306 94102
rect 39374 94046 39430 94102
rect 39498 94046 39554 94102
rect 39622 94046 39678 94102
rect 39250 93922 39306 93978
rect 39374 93922 39430 93978
rect 39498 93922 39554 93978
rect 39622 93922 39678 93978
rect 39250 76294 39306 76350
rect 39374 76294 39430 76350
rect 39498 76294 39554 76350
rect 39622 76294 39678 76350
rect 39250 76170 39306 76226
rect 39374 76170 39430 76226
rect 39498 76170 39554 76226
rect 39622 76170 39678 76226
rect 39250 76046 39306 76102
rect 39374 76046 39430 76102
rect 39498 76046 39554 76102
rect 39622 76046 39678 76102
rect 39250 75922 39306 75978
rect 39374 75922 39430 75978
rect 39498 75922 39554 75978
rect 39622 75922 39678 75978
rect 39250 58294 39306 58350
rect 39374 58294 39430 58350
rect 39498 58294 39554 58350
rect 39622 58294 39678 58350
rect 39250 58170 39306 58226
rect 39374 58170 39430 58226
rect 39498 58170 39554 58226
rect 39622 58170 39678 58226
rect 39250 58046 39306 58102
rect 39374 58046 39430 58102
rect 39498 58046 39554 58102
rect 39622 58046 39678 58102
rect 39250 57922 39306 57978
rect 39374 57922 39430 57978
rect 39498 57922 39554 57978
rect 39622 57922 39678 57978
rect 39250 40294 39306 40350
rect 39374 40294 39430 40350
rect 39498 40294 39554 40350
rect 39622 40294 39678 40350
rect 39250 40170 39306 40226
rect 39374 40170 39430 40226
rect 39498 40170 39554 40226
rect 39622 40170 39678 40226
rect 39250 40046 39306 40102
rect 39374 40046 39430 40102
rect 39498 40046 39554 40102
rect 39622 40046 39678 40102
rect 39250 39922 39306 39978
rect 39374 39922 39430 39978
rect 39498 39922 39554 39978
rect 39622 39922 39678 39978
rect 39250 22294 39306 22350
rect 39374 22294 39430 22350
rect 39498 22294 39554 22350
rect 39622 22294 39678 22350
rect 39250 22170 39306 22226
rect 39374 22170 39430 22226
rect 39498 22170 39554 22226
rect 39622 22170 39678 22226
rect 39250 22046 39306 22102
rect 39374 22046 39430 22102
rect 39498 22046 39554 22102
rect 39622 22046 39678 22102
rect 39250 21922 39306 21978
rect 39374 21922 39430 21978
rect 39498 21922 39554 21978
rect 39622 21922 39678 21978
rect 39250 4294 39306 4350
rect 39374 4294 39430 4350
rect 39498 4294 39554 4350
rect 39622 4294 39678 4350
rect 39250 4170 39306 4226
rect 39374 4170 39430 4226
rect 39498 4170 39554 4226
rect 39622 4170 39678 4226
rect 39250 4046 39306 4102
rect 39374 4046 39430 4102
rect 39498 4046 39554 4102
rect 39622 4046 39678 4102
rect 39250 3922 39306 3978
rect 39374 3922 39430 3978
rect 39498 3922 39554 3978
rect 39622 3922 39678 3978
rect 39250 -216 39306 -160
rect 39374 -216 39430 -160
rect 39498 -216 39554 -160
rect 39622 -216 39678 -160
rect 39250 -340 39306 -284
rect 39374 -340 39430 -284
rect 39498 -340 39554 -284
rect 39622 -340 39678 -284
rect 39250 -464 39306 -408
rect 39374 -464 39430 -408
rect 39498 -464 39554 -408
rect 39622 -464 39678 -408
rect 39250 -588 39306 -532
rect 39374 -588 39430 -532
rect 39498 -588 39554 -532
rect 39622 -588 39678 -532
rect 42970 598116 43026 598172
rect 43094 598116 43150 598172
rect 43218 598116 43274 598172
rect 43342 598116 43398 598172
rect 42970 597992 43026 598048
rect 43094 597992 43150 598048
rect 43218 597992 43274 598048
rect 43342 597992 43398 598048
rect 42970 597868 43026 597924
rect 43094 597868 43150 597924
rect 43218 597868 43274 597924
rect 43342 597868 43398 597924
rect 42970 597744 43026 597800
rect 43094 597744 43150 597800
rect 43218 597744 43274 597800
rect 43342 597744 43398 597800
rect 42970 586294 43026 586350
rect 43094 586294 43150 586350
rect 43218 586294 43274 586350
rect 43342 586294 43398 586350
rect 42970 586170 43026 586226
rect 43094 586170 43150 586226
rect 43218 586170 43274 586226
rect 43342 586170 43398 586226
rect 42970 586046 43026 586102
rect 43094 586046 43150 586102
rect 43218 586046 43274 586102
rect 43342 586046 43398 586102
rect 42970 585922 43026 585978
rect 43094 585922 43150 585978
rect 43218 585922 43274 585978
rect 43342 585922 43398 585978
rect 42970 568294 43026 568350
rect 43094 568294 43150 568350
rect 43218 568294 43274 568350
rect 43342 568294 43398 568350
rect 42970 568170 43026 568226
rect 43094 568170 43150 568226
rect 43218 568170 43274 568226
rect 43342 568170 43398 568226
rect 42970 568046 43026 568102
rect 43094 568046 43150 568102
rect 43218 568046 43274 568102
rect 43342 568046 43398 568102
rect 42970 567922 43026 567978
rect 43094 567922 43150 567978
rect 43218 567922 43274 567978
rect 43342 567922 43398 567978
rect 42970 550294 43026 550350
rect 43094 550294 43150 550350
rect 43218 550294 43274 550350
rect 43342 550294 43398 550350
rect 42970 550170 43026 550226
rect 43094 550170 43150 550226
rect 43218 550170 43274 550226
rect 43342 550170 43398 550226
rect 42970 550046 43026 550102
rect 43094 550046 43150 550102
rect 43218 550046 43274 550102
rect 43342 550046 43398 550102
rect 42970 549922 43026 549978
rect 43094 549922 43150 549978
rect 43218 549922 43274 549978
rect 43342 549922 43398 549978
rect 42970 532294 43026 532350
rect 43094 532294 43150 532350
rect 43218 532294 43274 532350
rect 43342 532294 43398 532350
rect 42970 532170 43026 532226
rect 43094 532170 43150 532226
rect 43218 532170 43274 532226
rect 43342 532170 43398 532226
rect 42970 532046 43026 532102
rect 43094 532046 43150 532102
rect 43218 532046 43274 532102
rect 43342 532046 43398 532102
rect 42970 531922 43026 531978
rect 43094 531922 43150 531978
rect 43218 531922 43274 531978
rect 43342 531922 43398 531978
rect 57250 597156 57306 597212
rect 57374 597156 57430 597212
rect 57498 597156 57554 597212
rect 57622 597156 57678 597212
rect 57250 597032 57306 597088
rect 57374 597032 57430 597088
rect 57498 597032 57554 597088
rect 57622 597032 57678 597088
rect 57250 596908 57306 596964
rect 57374 596908 57430 596964
rect 57498 596908 57554 596964
rect 57622 596908 57678 596964
rect 57250 596784 57306 596840
rect 57374 596784 57430 596840
rect 57498 596784 57554 596840
rect 57622 596784 57678 596840
rect 57250 580294 57306 580350
rect 57374 580294 57430 580350
rect 57498 580294 57554 580350
rect 57622 580294 57678 580350
rect 57250 580170 57306 580226
rect 57374 580170 57430 580226
rect 57498 580170 57554 580226
rect 57622 580170 57678 580226
rect 57250 580046 57306 580102
rect 57374 580046 57430 580102
rect 57498 580046 57554 580102
rect 57622 580046 57678 580102
rect 57250 579922 57306 579978
rect 57374 579922 57430 579978
rect 57498 579922 57554 579978
rect 57622 579922 57678 579978
rect 57250 562294 57306 562350
rect 57374 562294 57430 562350
rect 57498 562294 57554 562350
rect 57622 562294 57678 562350
rect 57250 562170 57306 562226
rect 57374 562170 57430 562226
rect 57498 562170 57554 562226
rect 57622 562170 57678 562226
rect 57250 562046 57306 562102
rect 57374 562046 57430 562102
rect 57498 562046 57554 562102
rect 57622 562046 57678 562102
rect 57250 561922 57306 561978
rect 57374 561922 57430 561978
rect 57498 561922 57554 561978
rect 57622 561922 57678 561978
rect 57250 544294 57306 544350
rect 57374 544294 57430 544350
rect 57498 544294 57554 544350
rect 57622 544294 57678 544350
rect 57250 544170 57306 544226
rect 57374 544170 57430 544226
rect 57498 544170 57554 544226
rect 57622 544170 57678 544226
rect 57250 544046 57306 544102
rect 57374 544046 57430 544102
rect 57498 544046 57554 544102
rect 57622 544046 57678 544102
rect 57250 543922 57306 543978
rect 57374 543922 57430 543978
rect 57498 543922 57554 543978
rect 57622 543922 57678 543978
rect 54518 526237 54574 526293
rect 54642 526237 54698 526293
rect 54518 526113 54574 526169
rect 54642 526113 54698 526169
rect 54518 525989 54574 526045
rect 54642 525989 54698 526045
rect 54518 525865 54574 525921
rect 54642 525865 54698 525921
rect 57250 526294 57306 526350
rect 57374 526294 57430 526350
rect 57498 526294 57554 526350
rect 57622 526294 57678 526350
rect 57250 526170 57306 526226
rect 57374 526170 57430 526226
rect 57498 526170 57554 526226
rect 57622 526170 57678 526226
rect 57250 526046 57306 526102
rect 57374 526046 57430 526102
rect 57498 526046 57554 526102
rect 57622 526046 57678 526102
rect 57250 525922 57306 525978
rect 57374 525922 57430 525978
rect 57498 525922 57554 525978
rect 57622 525922 57678 525978
rect 42970 514294 43026 514350
rect 43094 514294 43150 514350
rect 43218 514294 43274 514350
rect 43342 514294 43398 514350
rect 42970 514170 43026 514226
rect 43094 514170 43150 514226
rect 43218 514170 43274 514226
rect 43342 514170 43398 514226
rect 42970 514046 43026 514102
rect 43094 514046 43150 514102
rect 43218 514046 43274 514102
rect 43342 514046 43398 514102
rect 42970 513922 43026 513978
rect 43094 513922 43150 513978
rect 43218 513922 43274 513978
rect 43342 513922 43398 513978
rect 54518 508294 54574 508350
rect 54642 508294 54698 508350
rect 54518 508170 54574 508226
rect 54642 508170 54698 508226
rect 54518 508046 54574 508102
rect 54642 508046 54698 508102
rect 54518 507922 54574 507978
rect 54642 507922 54698 507978
rect 57250 508294 57306 508350
rect 57374 508294 57430 508350
rect 57498 508294 57554 508350
rect 57622 508294 57678 508350
rect 57250 508170 57306 508226
rect 57374 508170 57430 508226
rect 57498 508170 57554 508226
rect 57622 508170 57678 508226
rect 57250 508046 57306 508102
rect 57374 508046 57430 508102
rect 57498 508046 57554 508102
rect 57622 508046 57678 508102
rect 57250 507922 57306 507978
rect 57374 507922 57430 507978
rect 57498 507922 57554 507978
rect 57622 507922 57678 507978
rect 42970 496294 43026 496350
rect 43094 496294 43150 496350
rect 43218 496294 43274 496350
rect 43342 496294 43398 496350
rect 42970 496170 43026 496226
rect 43094 496170 43150 496226
rect 43218 496170 43274 496226
rect 43342 496170 43398 496226
rect 42970 496046 43026 496102
rect 43094 496046 43150 496102
rect 43218 496046 43274 496102
rect 43342 496046 43398 496102
rect 42970 495922 43026 495978
rect 43094 495922 43150 495978
rect 43218 495922 43274 495978
rect 43342 495922 43398 495978
rect 54518 490294 54574 490350
rect 54642 490294 54698 490350
rect 54518 490170 54574 490226
rect 54642 490170 54698 490226
rect 54518 490046 54574 490102
rect 54642 490046 54698 490102
rect 54518 489922 54574 489978
rect 54642 489922 54698 489978
rect 57250 490294 57306 490350
rect 57374 490294 57430 490350
rect 57498 490294 57554 490350
rect 57622 490294 57678 490350
rect 57250 490170 57306 490226
rect 57374 490170 57430 490226
rect 57498 490170 57554 490226
rect 57622 490170 57678 490226
rect 57250 490046 57306 490102
rect 57374 490046 57430 490102
rect 57498 490046 57554 490102
rect 57622 490046 57678 490102
rect 57250 489922 57306 489978
rect 57374 489922 57430 489978
rect 57498 489922 57554 489978
rect 57622 489922 57678 489978
rect 42970 478294 43026 478350
rect 43094 478294 43150 478350
rect 43218 478294 43274 478350
rect 43342 478294 43398 478350
rect 42970 478170 43026 478226
rect 43094 478170 43150 478226
rect 43218 478170 43274 478226
rect 43342 478170 43398 478226
rect 42970 478046 43026 478102
rect 43094 478046 43150 478102
rect 43218 478046 43274 478102
rect 43342 478046 43398 478102
rect 42970 477922 43026 477978
rect 43094 477922 43150 477978
rect 43218 477922 43274 477978
rect 43342 477922 43398 477978
rect 54518 472294 54574 472350
rect 54642 472294 54698 472350
rect 54518 472170 54574 472226
rect 54642 472170 54698 472226
rect 54518 472046 54574 472102
rect 54642 472046 54698 472102
rect 54518 471922 54574 471978
rect 54642 471922 54698 471978
rect 57250 472294 57306 472350
rect 57374 472294 57430 472350
rect 57498 472294 57554 472350
rect 57622 472294 57678 472350
rect 57250 472170 57306 472226
rect 57374 472170 57430 472226
rect 57498 472170 57554 472226
rect 57622 472170 57678 472226
rect 57250 472046 57306 472102
rect 57374 472046 57430 472102
rect 57498 472046 57554 472102
rect 57622 472046 57678 472102
rect 57250 471922 57306 471978
rect 57374 471922 57430 471978
rect 57498 471922 57554 471978
rect 57622 471922 57678 471978
rect 42970 460294 43026 460350
rect 43094 460294 43150 460350
rect 43218 460294 43274 460350
rect 43342 460294 43398 460350
rect 42970 460170 43026 460226
rect 43094 460170 43150 460226
rect 43218 460170 43274 460226
rect 43342 460170 43398 460226
rect 42970 460046 43026 460102
rect 43094 460046 43150 460102
rect 43218 460046 43274 460102
rect 43342 460046 43398 460102
rect 42970 459922 43026 459978
rect 43094 459922 43150 459978
rect 43218 459922 43274 459978
rect 43342 459922 43398 459978
rect 54518 454294 54574 454350
rect 54642 454294 54698 454350
rect 54518 454170 54574 454226
rect 54642 454170 54698 454226
rect 54518 454046 54574 454102
rect 54642 454046 54698 454102
rect 54518 453922 54574 453978
rect 54642 453922 54698 453978
rect 57250 454294 57306 454350
rect 57374 454294 57430 454350
rect 57498 454294 57554 454350
rect 57622 454294 57678 454350
rect 57250 454170 57306 454226
rect 57374 454170 57430 454226
rect 57498 454170 57554 454226
rect 57622 454170 57678 454226
rect 57250 454046 57306 454102
rect 57374 454046 57430 454102
rect 57498 454046 57554 454102
rect 57622 454046 57678 454102
rect 57250 453922 57306 453978
rect 57374 453922 57430 453978
rect 57498 453922 57554 453978
rect 57622 453922 57678 453978
rect 42970 442294 43026 442350
rect 43094 442294 43150 442350
rect 43218 442294 43274 442350
rect 43342 442294 43398 442350
rect 42970 442170 43026 442226
rect 43094 442170 43150 442226
rect 43218 442170 43274 442226
rect 43342 442170 43398 442226
rect 42970 442046 43026 442102
rect 43094 442046 43150 442102
rect 43218 442046 43274 442102
rect 43342 442046 43398 442102
rect 42970 441922 43026 441978
rect 43094 441922 43150 441978
rect 43218 441922 43274 441978
rect 43342 441922 43398 441978
rect 54518 436294 54574 436350
rect 54642 436294 54698 436350
rect 54518 436170 54574 436226
rect 54642 436170 54698 436226
rect 54518 436046 54574 436102
rect 54642 436046 54698 436102
rect 54518 435922 54574 435978
rect 54642 435922 54698 435978
rect 57250 436294 57306 436350
rect 57374 436294 57430 436350
rect 57498 436294 57554 436350
rect 57622 436294 57678 436350
rect 57250 436170 57306 436226
rect 57374 436170 57430 436226
rect 57498 436170 57554 436226
rect 57622 436170 57678 436226
rect 57250 436046 57306 436102
rect 57374 436046 57430 436102
rect 57498 436046 57554 436102
rect 57622 436046 57678 436102
rect 57250 435922 57306 435978
rect 57374 435922 57430 435978
rect 57498 435922 57554 435978
rect 57622 435922 57678 435978
rect 42970 424294 43026 424350
rect 43094 424294 43150 424350
rect 43218 424294 43274 424350
rect 43342 424294 43398 424350
rect 42970 424170 43026 424226
rect 43094 424170 43150 424226
rect 43218 424170 43274 424226
rect 43342 424170 43398 424226
rect 42970 424046 43026 424102
rect 43094 424046 43150 424102
rect 43218 424046 43274 424102
rect 43342 424046 43398 424102
rect 42970 423922 43026 423978
rect 43094 423922 43150 423978
rect 43218 423922 43274 423978
rect 43342 423922 43398 423978
rect 54518 418294 54574 418350
rect 54642 418294 54698 418350
rect 54518 418170 54574 418226
rect 54642 418170 54698 418226
rect 54518 418046 54574 418102
rect 54642 418046 54698 418102
rect 54518 417922 54574 417978
rect 54642 417922 54698 417978
rect 57250 418294 57306 418350
rect 57374 418294 57430 418350
rect 57498 418294 57554 418350
rect 57622 418294 57678 418350
rect 57250 418170 57306 418226
rect 57374 418170 57430 418226
rect 57498 418170 57554 418226
rect 57622 418170 57678 418226
rect 57250 418046 57306 418102
rect 57374 418046 57430 418102
rect 57498 418046 57554 418102
rect 57622 418046 57678 418102
rect 57250 417922 57306 417978
rect 57374 417922 57430 417978
rect 57498 417922 57554 417978
rect 57622 417922 57678 417978
rect 42970 406294 43026 406350
rect 43094 406294 43150 406350
rect 43218 406294 43274 406350
rect 43342 406294 43398 406350
rect 42970 406170 43026 406226
rect 43094 406170 43150 406226
rect 43218 406170 43274 406226
rect 43342 406170 43398 406226
rect 42970 406046 43026 406102
rect 43094 406046 43150 406102
rect 43218 406046 43274 406102
rect 43342 406046 43398 406102
rect 42970 405922 43026 405978
rect 43094 405922 43150 405978
rect 43218 405922 43274 405978
rect 43342 405922 43398 405978
rect 54518 400294 54574 400350
rect 54642 400294 54698 400350
rect 54518 400170 54574 400226
rect 54642 400170 54698 400226
rect 54518 400046 54574 400102
rect 54642 400046 54698 400102
rect 54518 399922 54574 399978
rect 54642 399922 54698 399978
rect 57250 400294 57306 400350
rect 57374 400294 57430 400350
rect 57498 400294 57554 400350
rect 57622 400294 57678 400350
rect 57250 400170 57306 400226
rect 57374 400170 57430 400226
rect 57498 400170 57554 400226
rect 57622 400170 57678 400226
rect 57250 400046 57306 400102
rect 57374 400046 57430 400102
rect 57498 400046 57554 400102
rect 57622 400046 57678 400102
rect 57250 399922 57306 399978
rect 57374 399922 57430 399978
rect 57498 399922 57554 399978
rect 57622 399922 57678 399978
rect 42970 388294 43026 388350
rect 43094 388294 43150 388350
rect 43218 388294 43274 388350
rect 43342 388294 43398 388350
rect 42970 388170 43026 388226
rect 43094 388170 43150 388226
rect 43218 388170 43274 388226
rect 43342 388170 43398 388226
rect 42970 388046 43026 388102
rect 43094 388046 43150 388102
rect 43218 388046 43274 388102
rect 43342 388046 43398 388102
rect 42970 387922 43026 387978
rect 43094 387922 43150 387978
rect 43218 387922 43274 387978
rect 43342 387922 43398 387978
rect 54518 382294 54574 382350
rect 54642 382294 54698 382350
rect 54518 382170 54574 382226
rect 54642 382170 54698 382226
rect 54518 382046 54574 382102
rect 54642 382046 54698 382102
rect 54518 381922 54574 381978
rect 54642 381922 54698 381978
rect 57250 382294 57306 382350
rect 57374 382294 57430 382350
rect 57498 382294 57554 382350
rect 57622 382294 57678 382350
rect 57250 382170 57306 382226
rect 57374 382170 57430 382226
rect 57498 382170 57554 382226
rect 57622 382170 57678 382226
rect 57250 382046 57306 382102
rect 57374 382046 57430 382102
rect 57498 382046 57554 382102
rect 57622 382046 57678 382102
rect 57250 381922 57306 381978
rect 57374 381922 57430 381978
rect 57498 381922 57554 381978
rect 57622 381922 57678 381978
rect 42970 370294 43026 370350
rect 43094 370294 43150 370350
rect 43218 370294 43274 370350
rect 43342 370294 43398 370350
rect 42970 370170 43026 370226
rect 43094 370170 43150 370226
rect 43218 370170 43274 370226
rect 43342 370170 43398 370226
rect 42970 370046 43026 370102
rect 43094 370046 43150 370102
rect 43218 370046 43274 370102
rect 43342 370046 43398 370102
rect 42970 369922 43026 369978
rect 43094 369922 43150 369978
rect 43218 369922 43274 369978
rect 43342 369922 43398 369978
rect 54518 364294 54574 364350
rect 54642 364294 54698 364350
rect 54518 364170 54574 364226
rect 54642 364170 54698 364226
rect 54518 364046 54574 364102
rect 54642 364046 54698 364102
rect 54518 363922 54574 363978
rect 54642 363922 54698 363978
rect 57250 364294 57306 364350
rect 57374 364294 57430 364350
rect 57498 364294 57554 364350
rect 57622 364294 57678 364350
rect 57250 364170 57306 364226
rect 57374 364170 57430 364226
rect 57498 364170 57554 364226
rect 57622 364170 57678 364226
rect 57250 364046 57306 364102
rect 57374 364046 57430 364102
rect 57498 364046 57554 364102
rect 57622 364046 57678 364102
rect 57250 363922 57306 363978
rect 57374 363922 57430 363978
rect 57498 363922 57554 363978
rect 57622 363922 57678 363978
rect 42970 352294 43026 352350
rect 43094 352294 43150 352350
rect 43218 352294 43274 352350
rect 43342 352294 43398 352350
rect 42970 352170 43026 352226
rect 43094 352170 43150 352226
rect 43218 352170 43274 352226
rect 43342 352170 43398 352226
rect 42970 352046 43026 352102
rect 43094 352046 43150 352102
rect 43218 352046 43274 352102
rect 43342 352046 43398 352102
rect 42970 351922 43026 351978
rect 43094 351922 43150 351978
rect 43218 351922 43274 351978
rect 43342 351922 43398 351978
rect 54518 346294 54574 346350
rect 54642 346294 54698 346350
rect 54518 346170 54574 346226
rect 54642 346170 54698 346226
rect 54518 346046 54574 346102
rect 54642 346046 54698 346102
rect 54518 345922 54574 345978
rect 54642 345922 54698 345978
rect 57250 346294 57306 346350
rect 57374 346294 57430 346350
rect 57498 346294 57554 346350
rect 57622 346294 57678 346350
rect 57250 346170 57306 346226
rect 57374 346170 57430 346226
rect 57498 346170 57554 346226
rect 57622 346170 57678 346226
rect 57250 346046 57306 346102
rect 57374 346046 57430 346102
rect 57498 346046 57554 346102
rect 57622 346046 57678 346102
rect 57250 345922 57306 345978
rect 57374 345922 57430 345978
rect 57498 345922 57554 345978
rect 57622 345922 57678 345978
rect 42970 334294 43026 334350
rect 43094 334294 43150 334350
rect 43218 334294 43274 334350
rect 43342 334294 43398 334350
rect 42970 334170 43026 334226
rect 43094 334170 43150 334226
rect 43218 334170 43274 334226
rect 43342 334170 43398 334226
rect 42970 334046 43026 334102
rect 43094 334046 43150 334102
rect 43218 334046 43274 334102
rect 43342 334046 43398 334102
rect 42970 333922 43026 333978
rect 43094 333922 43150 333978
rect 43218 333922 43274 333978
rect 43342 333922 43398 333978
rect 54518 328294 54574 328350
rect 54642 328294 54698 328350
rect 54518 328170 54574 328226
rect 54642 328170 54698 328226
rect 54518 328046 54574 328102
rect 54642 328046 54698 328102
rect 54518 327922 54574 327978
rect 54642 327922 54698 327978
rect 57250 328294 57306 328350
rect 57374 328294 57430 328350
rect 57498 328294 57554 328350
rect 57622 328294 57678 328350
rect 57250 328170 57306 328226
rect 57374 328170 57430 328226
rect 57498 328170 57554 328226
rect 57622 328170 57678 328226
rect 57250 328046 57306 328102
rect 57374 328046 57430 328102
rect 57498 328046 57554 328102
rect 57622 328046 57678 328102
rect 57250 327922 57306 327978
rect 57374 327922 57430 327978
rect 57498 327922 57554 327978
rect 57622 327922 57678 327978
rect 42970 316294 43026 316350
rect 43094 316294 43150 316350
rect 43218 316294 43274 316350
rect 43342 316294 43398 316350
rect 42970 316170 43026 316226
rect 43094 316170 43150 316226
rect 43218 316170 43274 316226
rect 43342 316170 43398 316226
rect 42970 316046 43026 316102
rect 43094 316046 43150 316102
rect 43218 316046 43274 316102
rect 43342 316046 43398 316102
rect 42970 315922 43026 315978
rect 43094 315922 43150 315978
rect 43218 315922 43274 315978
rect 43342 315922 43398 315978
rect 54518 310294 54574 310350
rect 54642 310294 54698 310350
rect 54518 310170 54574 310226
rect 54642 310170 54698 310226
rect 54518 310046 54574 310102
rect 54642 310046 54698 310102
rect 54518 309922 54574 309978
rect 54642 309922 54698 309978
rect 57250 310294 57306 310350
rect 57374 310294 57430 310350
rect 57498 310294 57554 310350
rect 57622 310294 57678 310350
rect 57250 310170 57306 310226
rect 57374 310170 57430 310226
rect 57498 310170 57554 310226
rect 57622 310170 57678 310226
rect 57250 310046 57306 310102
rect 57374 310046 57430 310102
rect 57498 310046 57554 310102
rect 57622 310046 57678 310102
rect 57250 309922 57306 309978
rect 57374 309922 57430 309978
rect 57498 309922 57554 309978
rect 57622 309922 57678 309978
rect 42970 298294 43026 298350
rect 43094 298294 43150 298350
rect 43218 298294 43274 298350
rect 43342 298294 43398 298350
rect 42970 298170 43026 298226
rect 43094 298170 43150 298226
rect 43218 298170 43274 298226
rect 43342 298170 43398 298226
rect 42970 298046 43026 298102
rect 43094 298046 43150 298102
rect 43218 298046 43274 298102
rect 43342 298046 43398 298102
rect 42970 297922 43026 297978
rect 43094 297922 43150 297978
rect 43218 297922 43274 297978
rect 43342 297922 43398 297978
rect 54518 292294 54574 292350
rect 54642 292294 54698 292350
rect 54518 292170 54574 292226
rect 54642 292170 54698 292226
rect 54518 292046 54574 292102
rect 54642 292046 54698 292102
rect 54518 291922 54574 291978
rect 54642 291922 54698 291978
rect 57250 292294 57306 292350
rect 57374 292294 57430 292350
rect 57498 292294 57554 292350
rect 57622 292294 57678 292350
rect 57250 292170 57306 292226
rect 57374 292170 57430 292226
rect 57498 292170 57554 292226
rect 57622 292170 57678 292226
rect 57250 292046 57306 292102
rect 57374 292046 57430 292102
rect 57498 292046 57554 292102
rect 57622 292046 57678 292102
rect 57250 291922 57306 291978
rect 57374 291922 57430 291978
rect 57498 291922 57554 291978
rect 57622 291922 57678 291978
rect 42970 280294 43026 280350
rect 43094 280294 43150 280350
rect 43218 280294 43274 280350
rect 43342 280294 43398 280350
rect 42970 280170 43026 280226
rect 43094 280170 43150 280226
rect 43218 280170 43274 280226
rect 43342 280170 43398 280226
rect 42970 280046 43026 280102
rect 43094 280046 43150 280102
rect 43218 280046 43274 280102
rect 43342 280046 43398 280102
rect 42970 279922 43026 279978
rect 43094 279922 43150 279978
rect 43218 279922 43274 279978
rect 43342 279922 43398 279978
rect 54518 274294 54574 274350
rect 54642 274294 54698 274350
rect 54518 274170 54574 274226
rect 54642 274170 54698 274226
rect 54518 274046 54574 274102
rect 54642 274046 54698 274102
rect 54518 273922 54574 273978
rect 54642 273922 54698 273978
rect 57250 274294 57306 274350
rect 57374 274294 57430 274350
rect 57498 274294 57554 274350
rect 57622 274294 57678 274350
rect 57250 274170 57306 274226
rect 57374 274170 57430 274226
rect 57498 274170 57554 274226
rect 57622 274170 57678 274226
rect 57250 274046 57306 274102
rect 57374 274046 57430 274102
rect 57498 274046 57554 274102
rect 57622 274046 57678 274102
rect 57250 273922 57306 273978
rect 57374 273922 57430 273978
rect 57498 273922 57554 273978
rect 57622 273922 57678 273978
rect 42970 262294 43026 262350
rect 43094 262294 43150 262350
rect 43218 262294 43274 262350
rect 43342 262294 43398 262350
rect 42970 262170 43026 262226
rect 43094 262170 43150 262226
rect 43218 262170 43274 262226
rect 43342 262170 43398 262226
rect 42970 262046 43026 262102
rect 43094 262046 43150 262102
rect 43218 262046 43274 262102
rect 43342 262046 43398 262102
rect 42970 261922 43026 261978
rect 43094 261922 43150 261978
rect 43218 261922 43274 261978
rect 43342 261922 43398 261978
rect 54518 256294 54574 256350
rect 54642 256294 54698 256350
rect 54518 256170 54574 256226
rect 54642 256170 54698 256226
rect 54518 256046 54574 256102
rect 54642 256046 54698 256102
rect 54518 255922 54574 255978
rect 54642 255922 54698 255978
rect 57250 256294 57306 256350
rect 57374 256294 57430 256350
rect 57498 256294 57554 256350
rect 57622 256294 57678 256350
rect 57250 256170 57306 256226
rect 57374 256170 57430 256226
rect 57498 256170 57554 256226
rect 57622 256170 57678 256226
rect 57250 256046 57306 256102
rect 57374 256046 57430 256102
rect 57498 256046 57554 256102
rect 57622 256046 57678 256102
rect 57250 255922 57306 255978
rect 57374 255922 57430 255978
rect 57498 255922 57554 255978
rect 57622 255922 57678 255978
rect 42970 244294 43026 244350
rect 43094 244294 43150 244350
rect 43218 244294 43274 244350
rect 43342 244294 43398 244350
rect 42970 244170 43026 244226
rect 43094 244170 43150 244226
rect 43218 244170 43274 244226
rect 43342 244170 43398 244226
rect 42970 244046 43026 244102
rect 43094 244046 43150 244102
rect 43218 244046 43274 244102
rect 43342 244046 43398 244102
rect 42970 243922 43026 243978
rect 43094 243922 43150 243978
rect 43218 243922 43274 243978
rect 43342 243922 43398 243978
rect 54518 238294 54574 238350
rect 54642 238294 54698 238350
rect 54518 238170 54574 238226
rect 54642 238170 54698 238226
rect 54518 238046 54574 238102
rect 54642 238046 54698 238102
rect 54518 237922 54574 237978
rect 54642 237922 54698 237978
rect 57250 238294 57306 238350
rect 57374 238294 57430 238350
rect 57498 238294 57554 238350
rect 57622 238294 57678 238350
rect 57250 238170 57306 238226
rect 57374 238170 57430 238226
rect 57498 238170 57554 238226
rect 57622 238170 57678 238226
rect 57250 238046 57306 238102
rect 57374 238046 57430 238102
rect 57498 238046 57554 238102
rect 57622 238046 57678 238102
rect 57250 237922 57306 237978
rect 57374 237922 57430 237978
rect 57498 237922 57554 237978
rect 57622 237922 57678 237978
rect 42970 226294 43026 226350
rect 43094 226294 43150 226350
rect 43218 226294 43274 226350
rect 43342 226294 43398 226350
rect 42970 226170 43026 226226
rect 43094 226170 43150 226226
rect 43218 226170 43274 226226
rect 43342 226170 43398 226226
rect 42970 226046 43026 226102
rect 43094 226046 43150 226102
rect 43218 226046 43274 226102
rect 43342 226046 43398 226102
rect 42970 225922 43026 225978
rect 43094 225922 43150 225978
rect 43218 225922 43274 225978
rect 43342 225922 43398 225978
rect 54518 220294 54574 220350
rect 54642 220294 54698 220350
rect 54518 220170 54574 220226
rect 54642 220170 54698 220226
rect 54518 220046 54574 220102
rect 54642 220046 54698 220102
rect 54518 219922 54574 219978
rect 54642 219922 54698 219978
rect 57250 220294 57306 220350
rect 57374 220294 57430 220350
rect 57498 220294 57554 220350
rect 57622 220294 57678 220350
rect 57250 220170 57306 220226
rect 57374 220170 57430 220226
rect 57498 220170 57554 220226
rect 57622 220170 57678 220226
rect 57250 220046 57306 220102
rect 57374 220046 57430 220102
rect 57498 220046 57554 220102
rect 57622 220046 57678 220102
rect 57250 219922 57306 219978
rect 57374 219922 57430 219978
rect 57498 219922 57554 219978
rect 57622 219922 57678 219978
rect 42970 208294 43026 208350
rect 43094 208294 43150 208350
rect 43218 208294 43274 208350
rect 43342 208294 43398 208350
rect 42970 208170 43026 208226
rect 43094 208170 43150 208226
rect 43218 208170 43274 208226
rect 43342 208170 43398 208226
rect 42970 208046 43026 208102
rect 43094 208046 43150 208102
rect 43218 208046 43274 208102
rect 43342 208046 43398 208102
rect 42970 207922 43026 207978
rect 43094 207922 43150 207978
rect 43218 207922 43274 207978
rect 43342 207922 43398 207978
rect 54518 202294 54574 202350
rect 54642 202294 54698 202350
rect 54518 202170 54574 202226
rect 54642 202170 54698 202226
rect 54518 202046 54574 202102
rect 54642 202046 54698 202102
rect 54518 201922 54574 201978
rect 54642 201922 54698 201978
rect 57250 202294 57306 202350
rect 57374 202294 57430 202350
rect 57498 202294 57554 202350
rect 57622 202294 57678 202350
rect 57250 202170 57306 202226
rect 57374 202170 57430 202226
rect 57498 202170 57554 202226
rect 57622 202170 57678 202226
rect 57250 202046 57306 202102
rect 57374 202046 57430 202102
rect 57498 202046 57554 202102
rect 57622 202046 57678 202102
rect 57250 201922 57306 201978
rect 57374 201922 57430 201978
rect 57498 201922 57554 201978
rect 57622 201922 57678 201978
rect 42970 190294 43026 190350
rect 43094 190294 43150 190350
rect 43218 190294 43274 190350
rect 43342 190294 43398 190350
rect 42970 190170 43026 190226
rect 43094 190170 43150 190226
rect 43218 190170 43274 190226
rect 43342 190170 43398 190226
rect 42970 190046 43026 190102
rect 43094 190046 43150 190102
rect 43218 190046 43274 190102
rect 43342 190046 43398 190102
rect 42970 189922 43026 189978
rect 43094 189922 43150 189978
rect 43218 189922 43274 189978
rect 43342 189922 43398 189978
rect 54518 184294 54574 184350
rect 54642 184294 54698 184350
rect 54518 184170 54574 184226
rect 54642 184170 54698 184226
rect 54518 184046 54574 184102
rect 54642 184046 54698 184102
rect 54518 183922 54574 183978
rect 54642 183922 54698 183978
rect 57250 184294 57306 184350
rect 57374 184294 57430 184350
rect 57498 184294 57554 184350
rect 57622 184294 57678 184350
rect 57250 184170 57306 184226
rect 57374 184170 57430 184226
rect 57498 184170 57554 184226
rect 57622 184170 57678 184226
rect 57250 184046 57306 184102
rect 57374 184046 57430 184102
rect 57498 184046 57554 184102
rect 57622 184046 57678 184102
rect 57250 183922 57306 183978
rect 57374 183922 57430 183978
rect 57498 183922 57554 183978
rect 57622 183922 57678 183978
rect 42970 172294 43026 172350
rect 43094 172294 43150 172350
rect 43218 172294 43274 172350
rect 43342 172294 43398 172350
rect 42970 172170 43026 172226
rect 43094 172170 43150 172226
rect 43218 172170 43274 172226
rect 43342 172170 43398 172226
rect 42970 172046 43026 172102
rect 43094 172046 43150 172102
rect 43218 172046 43274 172102
rect 43342 172046 43398 172102
rect 42970 171922 43026 171978
rect 43094 171922 43150 171978
rect 43218 171922 43274 171978
rect 43342 171922 43398 171978
rect 54518 166294 54574 166350
rect 54642 166294 54698 166350
rect 54518 166170 54574 166226
rect 54642 166170 54698 166226
rect 54518 166046 54574 166102
rect 54642 166046 54698 166102
rect 54518 165922 54574 165978
rect 54642 165922 54698 165978
rect 57250 166294 57306 166350
rect 57374 166294 57430 166350
rect 57498 166294 57554 166350
rect 57622 166294 57678 166350
rect 57250 166170 57306 166226
rect 57374 166170 57430 166226
rect 57498 166170 57554 166226
rect 57622 166170 57678 166226
rect 57250 166046 57306 166102
rect 57374 166046 57430 166102
rect 57498 166046 57554 166102
rect 57622 166046 57678 166102
rect 57250 165922 57306 165978
rect 57374 165922 57430 165978
rect 57498 165922 57554 165978
rect 57622 165922 57678 165978
rect 42970 154294 43026 154350
rect 43094 154294 43150 154350
rect 43218 154294 43274 154350
rect 43342 154294 43398 154350
rect 42970 154170 43026 154226
rect 43094 154170 43150 154226
rect 43218 154170 43274 154226
rect 43342 154170 43398 154226
rect 42970 154046 43026 154102
rect 43094 154046 43150 154102
rect 43218 154046 43274 154102
rect 43342 154046 43398 154102
rect 42970 153922 43026 153978
rect 43094 153922 43150 153978
rect 43218 153922 43274 153978
rect 43342 153922 43398 153978
rect 54518 148294 54574 148350
rect 54642 148294 54698 148350
rect 54518 148170 54574 148226
rect 54642 148170 54698 148226
rect 54518 148046 54574 148102
rect 54642 148046 54698 148102
rect 54518 147922 54574 147978
rect 54642 147922 54698 147978
rect 57250 148294 57306 148350
rect 57374 148294 57430 148350
rect 57498 148294 57554 148350
rect 57622 148294 57678 148350
rect 57250 148170 57306 148226
rect 57374 148170 57430 148226
rect 57498 148170 57554 148226
rect 57622 148170 57678 148226
rect 57250 148046 57306 148102
rect 57374 148046 57430 148102
rect 57498 148046 57554 148102
rect 57622 148046 57678 148102
rect 57250 147922 57306 147978
rect 57374 147922 57430 147978
rect 57498 147922 57554 147978
rect 57622 147922 57678 147978
rect 42970 136294 43026 136350
rect 43094 136294 43150 136350
rect 43218 136294 43274 136350
rect 43342 136294 43398 136350
rect 42970 136170 43026 136226
rect 43094 136170 43150 136226
rect 43218 136170 43274 136226
rect 43342 136170 43398 136226
rect 42970 136046 43026 136102
rect 43094 136046 43150 136102
rect 43218 136046 43274 136102
rect 43342 136046 43398 136102
rect 42970 135922 43026 135978
rect 43094 135922 43150 135978
rect 43218 135922 43274 135978
rect 43342 135922 43398 135978
rect 54518 130294 54574 130350
rect 54642 130294 54698 130350
rect 54518 130170 54574 130226
rect 54642 130170 54698 130226
rect 54518 130046 54574 130102
rect 54642 130046 54698 130102
rect 54518 129922 54574 129978
rect 54642 129922 54698 129978
rect 57250 130294 57306 130350
rect 57374 130294 57430 130350
rect 57498 130294 57554 130350
rect 57622 130294 57678 130350
rect 57250 130170 57306 130226
rect 57374 130170 57430 130226
rect 57498 130170 57554 130226
rect 57622 130170 57678 130226
rect 57250 130046 57306 130102
rect 57374 130046 57430 130102
rect 57498 130046 57554 130102
rect 57622 130046 57678 130102
rect 57250 129922 57306 129978
rect 57374 129922 57430 129978
rect 57498 129922 57554 129978
rect 57622 129922 57678 129978
rect 42970 118294 43026 118350
rect 43094 118294 43150 118350
rect 43218 118294 43274 118350
rect 43342 118294 43398 118350
rect 42970 118170 43026 118226
rect 43094 118170 43150 118226
rect 43218 118170 43274 118226
rect 43342 118170 43398 118226
rect 42970 118046 43026 118102
rect 43094 118046 43150 118102
rect 43218 118046 43274 118102
rect 43342 118046 43398 118102
rect 42970 117922 43026 117978
rect 43094 117922 43150 117978
rect 43218 117922 43274 117978
rect 43342 117922 43398 117978
rect 54518 112294 54574 112350
rect 54642 112294 54698 112350
rect 54518 112170 54574 112226
rect 54642 112170 54698 112226
rect 54518 112046 54574 112102
rect 54642 112046 54698 112102
rect 54518 111922 54574 111978
rect 54642 111922 54698 111978
rect 57250 112294 57306 112350
rect 57374 112294 57430 112350
rect 57498 112294 57554 112350
rect 57622 112294 57678 112350
rect 57250 112170 57306 112226
rect 57374 112170 57430 112226
rect 57498 112170 57554 112226
rect 57622 112170 57678 112226
rect 57250 112046 57306 112102
rect 57374 112046 57430 112102
rect 57498 112046 57554 112102
rect 57622 112046 57678 112102
rect 57250 111922 57306 111978
rect 57374 111922 57430 111978
rect 57498 111922 57554 111978
rect 57622 111922 57678 111978
rect 42970 100294 43026 100350
rect 43094 100294 43150 100350
rect 43218 100294 43274 100350
rect 43342 100294 43398 100350
rect 42970 100170 43026 100226
rect 43094 100170 43150 100226
rect 43218 100170 43274 100226
rect 43342 100170 43398 100226
rect 42970 100046 43026 100102
rect 43094 100046 43150 100102
rect 43218 100046 43274 100102
rect 43342 100046 43398 100102
rect 42970 99922 43026 99978
rect 43094 99922 43150 99978
rect 43218 99922 43274 99978
rect 43342 99922 43398 99978
rect 54518 94294 54574 94350
rect 54642 94294 54698 94350
rect 54518 94170 54574 94226
rect 54642 94170 54698 94226
rect 54518 94046 54574 94102
rect 54642 94046 54698 94102
rect 54518 93922 54574 93978
rect 54642 93922 54698 93978
rect 57250 94294 57306 94350
rect 57374 94294 57430 94350
rect 57498 94294 57554 94350
rect 57622 94294 57678 94350
rect 57250 94170 57306 94226
rect 57374 94170 57430 94226
rect 57498 94170 57554 94226
rect 57622 94170 57678 94226
rect 57250 94046 57306 94102
rect 57374 94046 57430 94102
rect 57498 94046 57554 94102
rect 57622 94046 57678 94102
rect 57250 93922 57306 93978
rect 57374 93922 57430 93978
rect 57498 93922 57554 93978
rect 57622 93922 57678 93978
rect 42970 82294 43026 82350
rect 43094 82294 43150 82350
rect 43218 82294 43274 82350
rect 43342 82294 43398 82350
rect 42970 82170 43026 82226
rect 43094 82170 43150 82226
rect 43218 82170 43274 82226
rect 43342 82170 43398 82226
rect 42970 82046 43026 82102
rect 43094 82046 43150 82102
rect 43218 82046 43274 82102
rect 43342 82046 43398 82102
rect 42970 81922 43026 81978
rect 43094 81922 43150 81978
rect 43218 81922 43274 81978
rect 43342 81922 43398 81978
rect 54518 76294 54574 76350
rect 54642 76294 54698 76350
rect 54518 76170 54574 76226
rect 54642 76170 54698 76226
rect 54518 76046 54574 76102
rect 54642 76046 54698 76102
rect 54518 75922 54574 75978
rect 54642 75922 54698 75978
rect 57250 76294 57306 76350
rect 57374 76294 57430 76350
rect 57498 76294 57554 76350
rect 57622 76294 57678 76350
rect 57250 76170 57306 76226
rect 57374 76170 57430 76226
rect 57498 76170 57554 76226
rect 57622 76170 57678 76226
rect 57250 76046 57306 76102
rect 57374 76046 57430 76102
rect 57498 76046 57554 76102
rect 57622 76046 57678 76102
rect 57250 75922 57306 75978
rect 57374 75922 57430 75978
rect 57498 75922 57554 75978
rect 57622 75922 57678 75978
rect 42970 64294 43026 64350
rect 43094 64294 43150 64350
rect 43218 64294 43274 64350
rect 43342 64294 43398 64350
rect 42970 64170 43026 64226
rect 43094 64170 43150 64226
rect 43218 64170 43274 64226
rect 43342 64170 43398 64226
rect 42970 64046 43026 64102
rect 43094 64046 43150 64102
rect 43218 64046 43274 64102
rect 43342 64046 43398 64102
rect 42970 63922 43026 63978
rect 43094 63922 43150 63978
rect 43218 63922 43274 63978
rect 43342 63922 43398 63978
rect 54518 58294 54574 58350
rect 54642 58294 54698 58350
rect 54518 58170 54574 58226
rect 54642 58170 54698 58226
rect 54518 58046 54574 58102
rect 54642 58046 54698 58102
rect 54518 57922 54574 57978
rect 54642 57922 54698 57978
rect 57250 58294 57306 58350
rect 57374 58294 57430 58350
rect 57498 58294 57554 58350
rect 57622 58294 57678 58350
rect 57250 58170 57306 58226
rect 57374 58170 57430 58226
rect 57498 58170 57554 58226
rect 57622 58170 57678 58226
rect 57250 58046 57306 58102
rect 57374 58046 57430 58102
rect 57498 58046 57554 58102
rect 57622 58046 57678 58102
rect 57250 57922 57306 57978
rect 57374 57922 57430 57978
rect 57498 57922 57554 57978
rect 57622 57922 57678 57978
rect 42970 46294 43026 46350
rect 43094 46294 43150 46350
rect 43218 46294 43274 46350
rect 43342 46294 43398 46350
rect 42970 46170 43026 46226
rect 43094 46170 43150 46226
rect 43218 46170 43274 46226
rect 43342 46170 43398 46226
rect 42970 46046 43026 46102
rect 43094 46046 43150 46102
rect 43218 46046 43274 46102
rect 43342 46046 43398 46102
rect 42970 45922 43026 45978
rect 43094 45922 43150 45978
rect 43218 45922 43274 45978
rect 43342 45922 43398 45978
rect 54518 40294 54574 40350
rect 54642 40294 54698 40350
rect 54518 40170 54574 40226
rect 54642 40170 54698 40226
rect 54518 40046 54574 40102
rect 54642 40046 54698 40102
rect 54518 39922 54574 39978
rect 54642 39922 54698 39978
rect 57250 40294 57306 40350
rect 57374 40294 57430 40350
rect 57498 40294 57554 40350
rect 57622 40294 57678 40350
rect 57250 40170 57306 40226
rect 57374 40170 57430 40226
rect 57498 40170 57554 40226
rect 57622 40170 57678 40226
rect 57250 40046 57306 40102
rect 57374 40046 57430 40102
rect 57498 40046 57554 40102
rect 57622 40046 57678 40102
rect 57250 39922 57306 39978
rect 57374 39922 57430 39978
rect 57498 39922 57554 39978
rect 57622 39922 57678 39978
rect 42970 28294 43026 28350
rect 43094 28294 43150 28350
rect 43218 28294 43274 28350
rect 43342 28294 43398 28350
rect 42970 28170 43026 28226
rect 43094 28170 43150 28226
rect 43218 28170 43274 28226
rect 43342 28170 43398 28226
rect 42970 28046 43026 28102
rect 43094 28046 43150 28102
rect 43218 28046 43274 28102
rect 43342 28046 43398 28102
rect 42970 27922 43026 27978
rect 43094 27922 43150 27978
rect 43218 27922 43274 27978
rect 43342 27922 43398 27978
rect 42970 10294 43026 10350
rect 43094 10294 43150 10350
rect 43218 10294 43274 10350
rect 43342 10294 43398 10350
rect 42970 10170 43026 10226
rect 43094 10170 43150 10226
rect 43218 10170 43274 10226
rect 43342 10170 43398 10226
rect 42970 10046 43026 10102
rect 43094 10046 43150 10102
rect 43218 10046 43274 10102
rect 43342 10046 43398 10102
rect 42970 9922 43026 9978
rect 43094 9922 43150 9978
rect 43218 9922 43274 9978
rect 43342 9922 43398 9978
rect 42970 -1176 43026 -1120
rect 43094 -1176 43150 -1120
rect 43218 -1176 43274 -1120
rect 43342 -1176 43398 -1120
rect 42970 -1300 43026 -1244
rect 43094 -1300 43150 -1244
rect 43218 -1300 43274 -1244
rect 43342 -1300 43398 -1244
rect 42970 -1424 43026 -1368
rect 43094 -1424 43150 -1368
rect 43218 -1424 43274 -1368
rect 43342 -1424 43398 -1368
rect 42970 -1548 43026 -1492
rect 43094 -1548 43150 -1492
rect 43218 -1548 43274 -1492
rect 43342 -1548 43398 -1492
rect 57250 22294 57306 22350
rect 57374 22294 57430 22350
rect 57498 22294 57554 22350
rect 57622 22294 57678 22350
rect 57250 22170 57306 22226
rect 57374 22170 57430 22226
rect 57498 22170 57554 22226
rect 57622 22170 57678 22226
rect 57250 22046 57306 22102
rect 57374 22046 57430 22102
rect 57498 22046 57554 22102
rect 57622 22046 57678 22102
rect 57250 21922 57306 21978
rect 57374 21922 57430 21978
rect 57498 21922 57554 21978
rect 57622 21922 57678 21978
rect 57250 4294 57306 4350
rect 57374 4294 57430 4350
rect 57498 4294 57554 4350
rect 57622 4294 57678 4350
rect 57250 4170 57306 4226
rect 57374 4170 57430 4226
rect 57498 4170 57554 4226
rect 57622 4170 57678 4226
rect 57250 4046 57306 4102
rect 57374 4046 57430 4102
rect 57498 4046 57554 4102
rect 57622 4046 57678 4102
rect 57250 3922 57306 3978
rect 57374 3922 57430 3978
rect 57498 3922 57554 3978
rect 57622 3922 57678 3978
rect 57250 -216 57306 -160
rect 57374 -216 57430 -160
rect 57498 -216 57554 -160
rect 57622 -216 57678 -160
rect 57250 -340 57306 -284
rect 57374 -340 57430 -284
rect 57498 -340 57554 -284
rect 57622 -340 57678 -284
rect 57250 -464 57306 -408
rect 57374 -464 57430 -408
rect 57498 -464 57554 -408
rect 57622 -464 57678 -408
rect 57250 -588 57306 -532
rect 57374 -588 57430 -532
rect 57498 -588 57554 -532
rect 57622 -588 57678 -532
rect 60970 598116 61026 598172
rect 61094 598116 61150 598172
rect 61218 598116 61274 598172
rect 61342 598116 61398 598172
rect 60970 597992 61026 598048
rect 61094 597992 61150 598048
rect 61218 597992 61274 598048
rect 61342 597992 61398 598048
rect 60970 597868 61026 597924
rect 61094 597868 61150 597924
rect 61218 597868 61274 597924
rect 61342 597868 61398 597924
rect 60970 597744 61026 597800
rect 61094 597744 61150 597800
rect 61218 597744 61274 597800
rect 61342 597744 61398 597800
rect 60970 586294 61026 586350
rect 61094 586294 61150 586350
rect 61218 586294 61274 586350
rect 61342 586294 61398 586350
rect 60970 586170 61026 586226
rect 61094 586170 61150 586226
rect 61218 586170 61274 586226
rect 61342 586170 61398 586226
rect 60970 586046 61026 586102
rect 61094 586046 61150 586102
rect 61218 586046 61274 586102
rect 61342 586046 61398 586102
rect 60970 585922 61026 585978
rect 61094 585922 61150 585978
rect 61218 585922 61274 585978
rect 61342 585922 61398 585978
rect 60970 568294 61026 568350
rect 61094 568294 61150 568350
rect 61218 568294 61274 568350
rect 61342 568294 61398 568350
rect 60970 568170 61026 568226
rect 61094 568170 61150 568226
rect 61218 568170 61274 568226
rect 61342 568170 61398 568226
rect 60970 568046 61026 568102
rect 61094 568046 61150 568102
rect 61218 568046 61274 568102
rect 61342 568046 61398 568102
rect 60970 567922 61026 567978
rect 61094 567922 61150 567978
rect 61218 567922 61274 567978
rect 61342 567922 61398 567978
rect 60970 550294 61026 550350
rect 61094 550294 61150 550350
rect 61218 550294 61274 550350
rect 61342 550294 61398 550350
rect 60970 550170 61026 550226
rect 61094 550170 61150 550226
rect 61218 550170 61274 550226
rect 61342 550170 61398 550226
rect 60970 550046 61026 550102
rect 61094 550046 61150 550102
rect 61218 550046 61274 550102
rect 61342 550046 61398 550102
rect 60970 549922 61026 549978
rect 61094 549922 61150 549978
rect 61218 549922 61274 549978
rect 61342 549922 61398 549978
rect 60970 532294 61026 532350
rect 61094 532294 61150 532350
rect 61218 532294 61274 532350
rect 61342 532294 61398 532350
rect 60970 532170 61026 532226
rect 61094 532170 61150 532226
rect 61218 532170 61274 532226
rect 61342 532170 61398 532226
rect 60970 532046 61026 532102
rect 61094 532046 61150 532102
rect 61218 532046 61274 532102
rect 61342 532046 61398 532102
rect 60970 531922 61026 531978
rect 61094 531922 61150 531978
rect 61218 531922 61274 531978
rect 61342 531922 61398 531978
rect 75250 597156 75306 597212
rect 75374 597156 75430 597212
rect 75498 597156 75554 597212
rect 75622 597156 75678 597212
rect 75250 597032 75306 597088
rect 75374 597032 75430 597088
rect 75498 597032 75554 597088
rect 75622 597032 75678 597088
rect 75250 596908 75306 596964
rect 75374 596908 75430 596964
rect 75498 596908 75554 596964
rect 75622 596908 75678 596964
rect 75250 596784 75306 596840
rect 75374 596784 75430 596840
rect 75498 596784 75554 596840
rect 75622 596784 75678 596840
rect 75250 580294 75306 580350
rect 75374 580294 75430 580350
rect 75498 580294 75554 580350
rect 75622 580294 75678 580350
rect 75250 580170 75306 580226
rect 75374 580170 75430 580226
rect 75498 580170 75554 580226
rect 75622 580170 75678 580226
rect 75250 580046 75306 580102
rect 75374 580046 75430 580102
rect 75498 580046 75554 580102
rect 75622 580046 75678 580102
rect 75250 579922 75306 579978
rect 75374 579922 75430 579978
rect 75498 579922 75554 579978
rect 75622 579922 75678 579978
rect 75250 562294 75306 562350
rect 75374 562294 75430 562350
rect 75498 562294 75554 562350
rect 75622 562294 75678 562350
rect 75250 562170 75306 562226
rect 75374 562170 75430 562226
rect 75498 562170 75554 562226
rect 75622 562170 75678 562226
rect 75250 562046 75306 562102
rect 75374 562046 75430 562102
rect 75498 562046 75554 562102
rect 75622 562046 75678 562102
rect 75250 561922 75306 561978
rect 75374 561922 75430 561978
rect 75498 561922 75554 561978
rect 75622 561922 75678 561978
rect 75250 544294 75306 544350
rect 75374 544294 75430 544350
rect 75498 544294 75554 544350
rect 75622 544294 75678 544350
rect 75250 544170 75306 544226
rect 75374 544170 75430 544226
rect 75498 544170 75554 544226
rect 75622 544170 75678 544226
rect 75250 544046 75306 544102
rect 75374 544046 75430 544102
rect 75498 544046 75554 544102
rect 75622 544046 75678 544102
rect 75250 543922 75306 543978
rect 75374 543922 75430 543978
rect 75498 543922 75554 543978
rect 75622 543922 75678 543978
rect 75250 526294 75306 526350
rect 75374 526294 75430 526350
rect 75498 526294 75554 526350
rect 75622 526294 75678 526350
rect 75250 526170 75306 526226
rect 75374 526170 75430 526226
rect 75498 526170 75554 526226
rect 75622 526170 75678 526226
rect 75250 526046 75306 526102
rect 75374 526046 75430 526102
rect 75498 526046 75554 526102
rect 75622 526046 75678 526102
rect 75250 525922 75306 525978
rect 75374 525922 75430 525978
rect 75498 525922 75554 525978
rect 75622 525922 75678 525978
rect 60970 514294 61026 514350
rect 61094 514294 61150 514350
rect 61218 514294 61274 514350
rect 61342 514294 61398 514350
rect 60970 514170 61026 514226
rect 61094 514170 61150 514226
rect 61218 514170 61274 514226
rect 61342 514170 61398 514226
rect 60970 514046 61026 514102
rect 61094 514046 61150 514102
rect 61218 514046 61274 514102
rect 61342 514046 61398 514102
rect 60970 513922 61026 513978
rect 61094 513922 61150 513978
rect 61218 513922 61274 513978
rect 61342 513922 61398 513978
rect 69878 514294 69934 514350
rect 70002 514294 70058 514350
rect 69878 514170 69934 514226
rect 70002 514170 70058 514226
rect 69878 514046 69934 514102
rect 70002 514046 70058 514102
rect 69878 513922 69934 513978
rect 70002 513922 70058 513978
rect 75250 508294 75306 508350
rect 75374 508294 75430 508350
rect 75498 508294 75554 508350
rect 75622 508294 75678 508350
rect 75250 508170 75306 508226
rect 75374 508170 75430 508226
rect 75498 508170 75554 508226
rect 75622 508170 75678 508226
rect 75250 508046 75306 508102
rect 75374 508046 75430 508102
rect 75498 508046 75554 508102
rect 75622 508046 75678 508102
rect 75250 507922 75306 507978
rect 75374 507922 75430 507978
rect 75498 507922 75554 507978
rect 75622 507922 75678 507978
rect 60970 496294 61026 496350
rect 61094 496294 61150 496350
rect 61218 496294 61274 496350
rect 61342 496294 61398 496350
rect 60970 496170 61026 496226
rect 61094 496170 61150 496226
rect 61218 496170 61274 496226
rect 61342 496170 61398 496226
rect 60970 496046 61026 496102
rect 61094 496046 61150 496102
rect 61218 496046 61274 496102
rect 61342 496046 61398 496102
rect 60970 495922 61026 495978
rect 61094 495922 61150 495978
rect 61218 495922 61274 495978
rect 61342 495922 61398 495978
rect 69878 496294 69934 496350
rect 70002 496294 70058 496350
rect 69878 496170 69934 496226
rect 70002 496170 70058 496226
rect 69878 496046 69934 496102
rect 70002 496046 70058 496102
rect 69878 495922 69934 495978
rect 70002 495922 70058 495978
rect 75250 490294 75306 490350
rect 75374 490294 75430 490350
rect 75498 490294 75554 490350
rect 75622 490294 75678 490350
rect 75250 490170 75306 490226
rect 75374 490170 75430 490226
rect 75498 490170 75554 490226
rect 75622 490170 75678 490226
rect 75250 490046 75306 490102
rect 75374 490046 75430 490102
rect 75498 490046 75554 490102
rect 75622 490046 75678 490102
rect 75250 489922 75306 489978
rect 75374 489922 75430 489978
rect 75498 489922 75554 489978
rect 75622 489922 75678 489978
rect 60970 478294 61026 478350
rect 61094 478294 61150 478350
rect 61218 478294 61274 478350
rect 61342 478294 61398 478350
rect 60970 478170 61026 478226
rect 61094 478170 61150 478226
rect 61218 478170 61274 478226
rect 61342 478170 61398 478226
rect 60970 478046 61026 478102
rect 61094 478046 61150 478102
rect 61218 478046 61274 478102
rect 61342 478046 61398 478102
rect 60970 477922 61026 477978
rect 61094 477922 61150 477978
rect 61218 477922 61274 477978
rect 61342 477922 61398 477978
rect 69878 478294 69934 478350
rect 70002 478294 70058 478350
rect 69878 478170 69934 478226
rect 70002 478170 70058 478226
rect 69878 478046 69934 478102
rect 70002 478046 70058 478102
rect 69878 477922 69934 477978
rect 70002 477922 70058 477978
rect 75250 472294 75306 472350
rect 75374 472294 75430 472350
rect 75498 472294 75554 472350
rect 75622 472294 75678 472350
rect 75250 472170 75306 472226
rect 75374 472170 75430 472226
rect 75498 472170 75554 472226
rect 75622 472170 75678 472226
rect 75250 472046 75306 472102
rect 75374 472046 75430 472102
rect 75498 472046 75554 472102
rect 75622 472046 75678 472102
rect 75250 471922 75306 471978
rect 75374 471922 75430 471978
rect 75498 471922 75554 471978
rect 75622 471922 75678 471978
rect 60970 460294 61026 460350
rect 61094 460294 61150 460350
rect 61218 460294 61274 460350
rect 61342 460294 61398 460350
rect 60970 460170 61026 460226
rect 61094 460170 61150 460226
rect 61218 460170 61274 460226
rect 61342 460170 61398 460226
rect 60970 460046 61026 460102
rect 61094 460046 61150 460102
rect 61218 460046 61274 460102
rect 61342 460046 61398 460102
rect 60970 459922 61026 459978
rect 61094 459922 61150 459978
rect 61218 459922 61274 459978
rect 61342 459922 61398 459978
rect 69878 460294 69934 460350
rect 70002 460294 70058 460350
rect 69878 460170 69934 460226
rect 70002 460170 70058 460226
rect 69878 460046 69934 460102
rect 70002 460046 70058 460102
rect 69878 459922 69934 459978
rect 70002 459922 70058 459978
rect 75250 454294 75306 454350
rect 75374 454294 75430 454350
rect 75498 454294 75554 454350
rect 75622 454294 75678 454350
rect 75250 454170 75306 454226
rect 75374 454170 75430 454226
rect 75498 454170 75554 454226
rect 75622 454170 75678 454226
rect 75250 454046 75306 454102
rect 75374 454046 75430 454102
rect 75498 454046 75554 454102
rect 75622 454046 75678 454102
rect 75250 453922 75306 453978
rect 75374 453922 75430 453978
rect 75498 453922 75554 453978
rect 75622 453922 75678 453978
rect 60970 442294 61026 442350
rect 61094 442294 61150 442350
rect 61218 442294 61274 442350
rect 61342 442294 61398 442350
rect 60970 442170 61026 442226
rect 61094 442170 61150 442226
rect 61218 442170 61274 442226
rect 61342 442170 61398 442226
rect 60970 442046 61026 442102
rect 61094 442046 61150 442102
rect 61218 442046 61274 442102
rect 61342 442046 61398 442102
rect 60970 441922 61026 441978
rect 61094 441922 61150 441978
rect 61218 441922 61274 441978
rect 61342 441922 61398 441978
rect 69878 442294 69934 442350
rect 70002 442294 70058 442350
rect 69878 442170 69934 442226
rect 70002 442170 70058 442226
rect 69878 442046 69934 442102
rect 70002 442046 70058 442102
rect 69878 441922 69934 441978
rect 70002 441922 70058 441978
rect 75250 436294 75306 436350
rect 75374 436294 75430 436350
rect 75498 436294 75554 436350
rect 75622 436294 75678 436350
rect 75250 436170 75306 436226
rect 75374 436170 75430 436226
rect 75498 436170 75554 436226
rect 75622 436170 75678 436226
rect 75250 436046 75306 436102
rect 75374 436046 75430 436102
rect 75498 436046 75554 436102
rect 75622 436046 75678 436102
rect 75250 435922 75306 435978
rect 75374 435922 75430 435978
rect 75498 435922 75554 435978
rect 75622 435922 75678 435978
rect 60970 424294 61026 424350
rect 61094 424294 61150 424350
rect 61218 424294 61274 424350
rect 61342 424294 61398 424350
rect 60970 424170 61026 424226
rect 61094 424170 61150 424226
rect 61218 424170 61274 424226
rect 61342 424170 61398 424226
rect 60970 424046 61026 424102
rect 61094 424046 61150 424102
rect 61218 424046 61274 424102
rect 61342 424046 61398 424102
rect 60970 423922 61026 423978
rect 61094 423922 61150 423978
rect 61218 423922 61274 423978
rect 61342 423922 61398 423978
rect 69878 424294 69934 424350
rect 70002 424294 70058 424350
rect 69878 424170 69934 424226
rect 70002 424170 70058 424226
rect 69878 424046 69934 424102
rect 70002 424046 70058 424102
rect 69878 423922 69934 423978
rect 70002 423922 70058 423978
rect 75250 418294 75306 418350
rect 75374 418294 75430 418350
rect 75498 418294 75554 418350
rect 75622 418294 75678 418350
rect 75250 418170 75306 418226
rect 75374 418170 75430 418226
rect 75498 418170 75554 418226
rect 75622 418170 75678 418226
rect 75250 418046 75306 418102
rect 75374 418046 75430 418102
rect 75498 418046 75554 418102
rect 75622 418046 75678 418102
rect 75250 417922 75306 417978
rect 75374 417922 75430 417978
rect 75498 417922 75554 417978
rect 75622 417922 75678 417978
rect 60970 406294 61026 406350
rect 61094 406294 61150 406350
rect 61218 406294 61274 406350
rect 61342 406294 61398 406350
rect 60970 406170 61026 406226
rect 61094 406170 61150 406226
rect 61218 406170 61274 406226
rect 61342 406170 61398 406226
rect 60970 406046 61026 406102
rect 61094 406046 61150 406102
rect 61218 406046 61274 406102
rect 61342 406046 61398 406102
rect 60970 405922 61026 405978
rect 61094 405922 61150 405978
rect 61218 405922 61274 405978
rect 61342 405922 61398 405978
rect 69878 406294 69934 406350
rect 70002 406294 70058 406350
rect 69878 406170 69934 406226
rect 70002 406170 70058 406226
rect 69878 406046 69934 406102
rect 70002 406046 70058 406102
rect 69878 405922 69934 405978
rect 70002 405922 70058 405978
rect 75250 400294 75306 400350
rect 75374 400294 75430 400350
rect 75498 400294 75554 400350
rect 75622 400294 75678 400350
rect 75250 400170 75306 400226
rect 75374 400170 75430 400226
rect 75498 400170 75554 400226
rect 75622 400170 75678 400226
rect 75250 400046 75306 400102
rect 75374 400046 75430 400102
rect 75498 400046 75554 400102
rect 75622 400046 75678 400102
rect 75250 399922 75306 399978
rect 75374 399922 75430 399978
rect 75498 399922 75554 399978
rect 75622 399922 75678 399978
rect 60970 388294 61026 388350
rect 61094 388294 61150 388350
rect 61218 388294 61274 388350
rect 61342 388294 61398 388350
rect 60970 388170 61026 388226
rect 61094 388170 61150 388226
rect 61218 388170 61274 388226
rect 61342 388170 61398 388226
rect 60970 388046 61026 388102
rect 61094 388046 61150 388102
rect 61218 388046 61274 388102
rect 61342 388046 61398 388102
rect 60970 387922 61026 387978
rect 61094 387922 61150 387978
rect 61218 387922 61274 387978
rect 61342 387922 61398 387978
rect 69878 388294 69934 388350
rect 70002 388294 70058 388350
rect 69878 388170 69934 388226
rect 70002 388170 70058 388226
rect 69878 388046 69934 388102
rect 70002 388046 70058 388102
rect 69878 387922 69934 387978
rect 70002 387922 70058 387978
rect 75250 382294 75306 382350
rect 75374 382294 75430 382350
rect 75498 382294 75554 382350
rect 75622 382294 75678 382350
rect 75250 382170 75306 382226
rect 75374 382170 75430 382226
rect 75498 382170 75554 382226
rect 75622 382170 75678 382226
rect 75250 382046 75306 382102
rect 75374 382046 75430 382102
rect 75498 382046 75554 382102
rect 75622 382046 75678 382102
rect 75250 381922 75306 381978
rect 75374 381922 75430 381978
rect 75498 381922 75554 381978
rect 75622 381922 75678 381978
rect 60970 370294 61026 370350
rect 61094 370294 61150 370350
rect 61218 370294 61274 370350
rect 61342 370294 61398 370350
rect 60970 370170 61026 370226
rect 61094 370170 61150 370226
rect 61218 370170 61274 370226
rect 61342 370170 61398 370226
rect 60970 370046 61026 370102
rect 61094 370046 61150 370102
rect 61218 370046 61274 370102
rect 61342 370046 61398 370102
rect 60970 369922 61026 369978
rect 61094 369922 61150 369978
rect 61218 369922 61274 369978
rect 61342 369922 61398 369978
rect 69878 370294 69934 370350
rect 70002 370294 70058 370350
rect 69878 370170 69934 370226
rect 70002 370170 70058 370226
rect 69878 370046 69934 370102
rect 70002 370046 70058 370102
rect 69878 369922 69934 369978
rect 70002 369922 70058 369978
rect 75250 364294 75306 364350
rect 75374 364294 75430 364350
rect 75498 364294 75554 364350
rect 75622 364294 75678 364350
rect 75250 364170 75306 364226
rect 75374 364170 75430 364226
rect 75498 364170 75554 364226
rect 75622 364170 75678 364226
rect 75250 364046 75306 364102
rect 75374 364046 75430 364102
rect 75498 364046 75554 364102
rect 75622 364046 75678 364102
rect 75250 363922 75306 363978
rect 75374 363922 75430 363978
rect 75498 363922 75554 363978
rect 75622 363922 75678 363978
rect 60970 352294 61026 352350
rect 61094 352294 61150 352350
rect 61218 352294 61274 352350
rect 61342 352294 61398 352350
rect 60970 352170 61026 352226
rect 61094 352170 61150 352226
rect 61218 352170 61274 352226
rect 61342 352170 61398 352226
rect 60970 352046 61026 352102
rect 61094 352046 61150 352102
rect 61218 352046 61274 352102
rect 61342 352046 61398 352102
rect 60970 351922 61026 351978
rect 61094 351922 61150 351978
rect 61218 351922 61274 351978
rect 61342 351922 61398 351978
rect 69878 352294 69934 352350
rect 70002 352294 70058 352350
rect 69878 352170 69934 352226
rect 70002 352170 70058 352226
rect 69878 352046 69934 352102
rect 70002 352046 70058 352102
rect 69878 351922 69934 351978
rect 70002 351922 70058 351978
rect 75250 346294 75306 346350
rect 75374 346294 75430 346350
rect 75498 346294 75554 346350
rect 75622 346294 75678 346350
rect 75250 346170 75306 346226
rect 75374 346170 75430 346226
rect 75498 346170 75554 346226
rect 75622 346170 75678 346226
rect 75250 346046 75306 346102
rect 75374 346046 75430 346102
rect 75498 346046 75554 346102
rect 75622 346046 75678 346102
rect 75250 345922 75306 345978
rect 75374 345922 75430 345978
rect 75498 345922 75554 345978
rect 75622 345922 75678 345978
rect 60970 334294 61026 334350
rect 61094 334294 61150 334350
rect 61218 334294 61274 334350
rect 61342 334294 61398 334350
rect 60970 334170 61026 334226
rect 61094 334170 61150 334226
rect 61218 334170 61274 334226
rect 61342 334170 61398 334226
rect 60970 334046 61026 334102
rect 61094 334046 61150 334102
rect 61218 334046 61274 334102
rect 61342 334046 61398 334102
rect 60970 333922 61026 333978
rect 61094 333922 61150 333978
rect 61218 333922 61274 333978
rect 61342 333922 61398 333978
rect 69878 334294 69934 334350
rect 70002 334294 70058 334350
rect 69878 334170 69934 334226
rect 70002 334170 70058 334226
rect 69878 334046 69934 334102
rect 70002 334046 70058 334102
rect 69878 333922 69934 333978
rect 70002 333922 70058 333978
rect 75250 328294 75306 328350
rect 75374 328294 75430 328350
rect 75498 328294 75554 328350
rect 75622 328294 75678 328350
rect 75250 328170 75306 328226
rect 75374 328170 75430 328226
rect 75498 328170 75554 328226
rect 75622 328170 75678 328226
rect 75250 328046 75306 328102
rect 75374 328046 75430 328102
rect 75498 328046 75554 328102
rect 75622 328046 75678 328102
rect 75250 327922 75306 327978
rect 75374 327922 75430 327978
rect 75498 327922 75554 327978
rect 75622 327922 75678 327978
rect 60970 316294 61026 316350
rect 61094 316294 61150 316350
rect 61218 316294 61274 316350
rect 61342 316294 61398 316350
rect 60970 316170 61026 316226
rect 61094 316170 61150 316226
rect 61218 316170 61274 316226
rect 61342 316170 61398 316226
rect 60970 316046 61026 316102
rect 61094 316046 61150 316102
rect 61218 316046 61274 316102
rect 61342 316046 61398 316102
rect 60970 315922 61026 315978
rect 61094 315922 61150 315978
rect 61218 315922 61274 315978
rect 61342 315922 61398 315978
rect 69878 316294 69934 316350
rect 70002 316294 70058 316350
rect 69878 316170 69934 316226
rect 70002 316170 70058 316226
rect 69878 316046 69934 316102
rect 70002 316046 70058 316102
rect 69878 315922 69934 315978
rect 70002 315922 70058 315978
rect 75250 310294 75306 310350
rect 75374 310294 75430 310350
rect 75498 310294 75554 310350
rect 75622 310294 75678 310350
rect 75250 310170 75306 310226
rect 75374 310170 75430 310226
rect 75498 310170 75554 310226
rect 75622 310170 75678 310226
rect 75250 310046 75306 310102
rect 75374 310046 75430 310102
rect 75498 310046 75554 310102
rect 75622 310046 75678 310102
rect 75250 309922 75306 309978
rect 75374 309922 75430 309978
rect 75498 309922 75554 309978
rect 75622 309922 75678 309978
rect 60970 298294 61026 298350
rect 61094 298294 61150 298350
rect 61218 298294 61274 298350
rect 61342 298294 61398 298350
rect 60970 298170 61026 298226
rect 61094 298170 61150 298226
rect 61218 298170 61274 298226
rect 61342 298170 61398 298226
rect 60970 298046 61026 298102
rect 61094 298046 61150 298102
rect 61218 298046 61274 298102
rect 61342 298046 61398 298102
rect 60970 297922 61026 297978
rect 61094 297922 61150 297978
rect 61218 297922 61274 297978
rect 61342 297922 61398 297978
rect 69878 298294 69934 298350
rect 70002 298294 70058 298350
rect 69878 298170 69934 298226
rect 70002 298170 70058 298226
rect 69878 298046 69934 298102
rect 70002 298046 70058 298102
rect 69878 297922 69934 297978
rect 70002 297922 70058 297978
rect 75250 292294 75306 292350
rect 75374 292294 75430 292350
rect 75498 292294 75554 292350
rect 75622 292294 75678 292350
rect 75250 292170 75306 292226
rect 75374 292170 75430 292226
rect 75498 292170 75554 292226
rect 75622 292170 75678 292226
rect 75250 292046 75306 292102
rect 75374 292046 75430 292102
rect 75498 292046 75554 292102
rect 75622 292046 75678 292102
rect 75250 291922 75306 291978
rect 75374 291922 75430 291978
rect 75498 291922 75554 291978
rect 75622 291922 75678 291978
rect 60970 280294 61026 280350
rect 61094 280294 61150 280350
rect 61218 280294 61274 280350
rect 61342 280294 61398 280350
rect 60970 280170 61026 280226
rect 61094 280170 61150 280226
rect 61218 280170 61274 280226
rect 61342 280170 61398 280226
rect 60970 280046 61026 280102
rect 61094 280046 61150 280102
rect 61218 280046 61274 280102
rect 61342 280046 61398 280102
rect 60970 279922 61026 279978
rect 61094 279922 61150 279978
rect 61218 279922 61274 279978
rect 61342 279922 61398 279978
rect 69878 280294 69934 280350
rect 70002 280294 70058 280350
rect 69878 280170 69934 280226
rect 70002 280170 70058 280226
rect 69878 280046 69934 280102
rect 70002 280046 70058 280102
rect 69878 279922 69934 279978
rect 70002 279922 70058 279978
rect 75250 274294 75306 274350
rect 75374 274294 75430 274350
rect 75498 274294 75554 274350
rect 75622 274294 75678 274350
rect 75250 274170 75306 274226
rect 75374 274170 75430 274226
rect 75498 274170 75554 274226
rect 75622 274170 75678 274226
rect 75250 274046 75306 274102
rect 75374 274046 75430 274102
rect 75498 274046 75554 274102
rect 75622 274046 75678 274102
rect 75250 273922 75306 273978
rect 75374 273922 75430 273978
rect 75498 273922 75554 273978
rect 75622 273922 75678 273978
rect 60970 262294 61026 262350
rect 61094 262294 61150 262350
rect 61218 262294 61274 262350
rect 61342 262294 61398 262350
rect 60970 262170 61026 262226
rect 61094 262170 61150 262226
rect 61218 262170 61274 262226
rect 61342 262170 61398 262226
rect 60970 262046 61026 262102
rect 61094 262046 61150 262102
rect 61218 262046 61274 262102
rect 61342 262046 61398 262102
rect 60970 261922 61026 261978
rect 61094 261922 61150 261978
rect 61218 261922 61274 261978
rect 61342 261922 61398 261978
rect 69878 262294 69934 262350
rect 70002 262294 70058 262350
rect 69878 262170 69934 262226
rect 70002 262170 70058 262226
rect 69878 262046 69934 262102
rect 70002 262046 70058 262102
rect 69878 261922 69934 261978
rect 70002 261922 70058 261978
rect 75250 256294 75306 256350
rect 75374 256294 75430 256350
rect 75498 256294 75554 256350
rect 75622 256294 75678 256350
rect 75250 256170 75306 256226
rect 75374 256170 75430 256226
rect 75498 256170 75554 256226
rect 75622 256170 75678 256226
rect 75250 256046 75306 256102
rect 75374 256046 75430 256102
rect 75498 256046 75554 256102
rect 75622 256046 75678 256102
rect 75250 255922 75306 255978
rect 75374 255922 75430 255978
rect 75498 255922 75554 255978
rect 75622 255922 75678 255978
rect 60970 244294 61026 244350
rect 61094 244294 61150 244350
rect 61218 244294 61274 244350
rect 61342 244294 61398 244350
rect 60970 244170 61026 244226
rect 61094 244170 61150 244226
rect 61218 244170 61274 244226
rect 61342 244170 61398 244226
rect 60970 244046 61026 244102
rect 61094 244046 61150 244102
rect 61218 244046 61274 244102
rect 61342 244046 61398 244102
rect 60970 243922 61026 243978
rect 61094 243922 61150 243978
rect 61218 243922 61274 243978
rect 61342 243922 61398 243978
rect 69878 244294 69934 244350
rect 70002 244294 70058 244350
rect 69878 244170 69934 244226
rect 70002 244170 70058 244226
rect 69878 244046 69934 244102
rect 70002 244046 70058 244102
rect 69878 243922 69934 243978
rect 70002 243922 70058 243978
rect 75250 238294 75306 238350
rect 75374 238294 75430 238350
rect 75498 238294 75554 238350
rect 75622 238294 75678 238350
rect 75250 238170 75306 238226
rect 75374 238170 75430 238226
rect 75498 238170 75554 238226
rect 75622 238170 75678 238226
rect 75250 238046 75306 238102
rect 75374 238046 75430 238102
rect 75498 238046 75554 238102
rect 75622 238046 75678 238102
rect 75250 237922 75306 237978
rect 75374 237922 75430 237978
rect 75498 237922 75554 237978
rect 75622 237922 75678 237978
rect 60970 226294 61026 226350
rect 61094 226294 61150 226350
rect 61218 226294 61274 226350
rect 61342 226294 61398 226350
rect 60970 226170 61026 226226
rect 61094 226170 61150 226226
rect 61218 226170 61274 226226
rect 61342 226170 61398 226226
rect 60970 226046 61026 226102
rect 61094 226046 61150 226102
rect 61218 226046 61274 226102
rect 61342 226046 61398 226102
rect 60970 225922 61026 225978
rect 61094 225922 61150 225978
rect 61218 225922 61274 225978
rect 61342 225922 61398 225978
rect 69878 226294 69934 226350
rect 70002 226294 70058 226350
rect 69878 226170 69934 226226
rect 70002 226170 70058 226226
rect 69878 226046 69934 226102
rect 70002 226046 70058 226102
rect 69878 225922 69934 225978
rect 70002 225922 70058 225978
rect 75250 220294 75306 220350
rect 75374 220294 75430 220350
rect 75498 220294 75554 220350
rect 75622 220294 75678 220350
rect 75250 220170 75306 220226
rect 75374 220170 75430 220226
rect 75498 220170 75554 220226
rect 75622 220170 75678 220226
rect 75250 220046 75306 220102
rect 75374 220046 75430 220102
rect 75498 220046 75554 220102
rect 75622 220046 75678 220102
rect 75250 219922 75306 219978
rect 75374 219922 75430 219978
rect 75498 219922 75554 219978
rect 75622 219922 75678 219978
rect 60970 208294 61026 208350
rect 61094 208294 61150 208350
rect 61218 208294 61274 208350
rect 61342 208294 61398 208350
rect 60970 208170 61026 208226
rect 61094 208170 61150 208226
rect 61218 208170 61274 208226
rect 61342 208170 61398 208226
rect 60970 208046 61026 208102
rect 61094 208046 61150 208102
rect 61218 208046 61274 208102
rect 61342 208046 61398 208102
rect 60970 207922 61026 207978
rect 61094 207922 61150 207978
rect 61218 207922 61274 207978
rect 61342 207922 61398 207978
rect 69878 208294 69934 208350
rect 70002 208294 70058 208350
rect 69878 208170 69934 208226
rect 70002 208170 70058 208226
rect 69878 208046 69934 208102
rect 70002 208046 70058 208102
rect 69878 207922 69934 207978
rect 70002 207922 70058 207978
rect 75250 202294 75306 202350
rect 75374 202294 75430 202350
rect 75498 202294 75554 202350
rect 75622 202294 75678 202350
rect 75250 202170 75306 202226
rect 75374 202170 75430 202226
rect 75498 202170 75554 202226
rect 75622 202170 75678 202226
rect 75250 202046 75306 202102
rect 75374 202046 75430 202102
rect 75498 202046 75554 202102
rect 75622 202046 75678 202102
rect 75250 201922 75306 201978
rect 75374 201922 75430 201978
rect 75498 201922 75554 201978
rect 75622 201922 75678 201978
rect 60970 190294 61026 190350
rect 61094 190294 61150 190350
rect 61218 190294 61274 190350
rect 61342 190294 61398 190350
rect 60970 190170 61026 190226
rect 61094 190170 61150 190226
rect 61218 190170 61274 190226
rect 61342 190170 61398 190226
rect 60970 190046 61026 190102
rect 61094 190046 61150 190102
rect 61218 190046 61274 190102
rect 61342 190046 61398 190102
rect 60970 189922 61026 189978
rect 61094 189922 61150 189978
rect 61218 189922 61274 189978
rect 61342 189922 61398 189978
rect 69878 190294 69934 190350
rect 70002 190294 70058 190350
rect 69878 190170 69934 190226
rect 70002 190170 70058 190226
rect 69878 190046 69934 190102
rect 70002 190046 70058 190102
rect 69878 189922 69934 189978
rect 70002 189922 70058 189978
rect 75250 184294 75306 184350
rect 75374 184294 75430 184350
rect 75498 184294 75554 184350
rect 75622 184294 75678 184350
rect 75250 184170 75306 184226
rect 75374 184170 75430 184226
rect 75498 184170 75554 184226
rect 75622 184170 75678 184226
rect 75250 184046 75306 184102
rect 75374 184046 75430 184102
rect 75498 184046 75554 184102
rect 75622 184046 75678 184102
rect 75250 183922 75306 183978
rect 75374 183922 75430 183978
rect 75498 183922 75554 183978
rect 75622 183922 75678 183978
rect 60970 172294 61026 172350
rect 61094 172294 61150 172350
rect 61218 172294 61274 172350
rect 61342 172294 61398 172350
rect 60970 172170 61026 172226
rect 61094 172170 61150 172226
rect 61218 172170 61274 172226
rect 61342 172170 61398 172226
rect 60970 172046 61026 172102
rect 61094 172046 61150 172102
rect 61218 172046 61274 172102
rect 61342 172046 61398 172102
rect 60970 171922 61026 171978
rect 61094 171922 61150 171978
rect 61218 171922 61274 171978
rect 61342 171922 61398 171978
rect 69878 172294 69934 172350
rect 70002 172294 70058 172350
rect 69878 172170 69934 172226
rect 70002 172170 70058 172226
rect 69878 172046 69934 172102
rect 70002 172046 70058 172102
rect 69878 171922 69934 171978
rect 70002 171922 70058 171978
rect 75250 166294 75306 166350
rect 75374 166294 75430 166350
rect 75498 166294 75554 166350
rect 75622 166294 75678 166350
rect 75250 166170 75306 166226
rect 75374 166170 75430 166226
rect 75498 166170 75554 166226
rect 75622 166170 75678 166226
rect 75250 166046 75306 166102
rect 75374 166046 75430 166102
rect 75498 166046 75554 166102
rect 75622 166046 75678 166102
rect 75250 165922 75306 165978
rect 75374 165922 75430 165978
rect 75498 165922 75554 165978
rect 75622 165922 75678 165978
rect 60970 154294 61026 154350
rect 61094 154294 61150 154350
rect 61218 154294 61274 154350
rect 61342 154294 61398 154350
rect 60970 154170 61026 154226
rect 61094 154170 61150 154226
rect 61218 154170 61274 154226
rect 61342 154170 61398 154226
rect 60970 154046 61026 154102
rect 61094 154046 61150 154102
rect 61218 154046 61274 154102
rect 61342 154046 61398 154102
rect 60970 153922 61026 153978
rect 61094 153922 61150 153978
rect 61218 153922 61274 153978
rect 61342 153922 61398 153978
rect 69878 154294 69934 154350
rect 70002 154294 70058 154350
rect 69878 154170 69934 154226
rect 70002 154170 70058 154226
rect 69878 154046 69934 154102
rect 70002 154046 70058 154102
rect 69878 153922 69934 153978
rect 70002 153922 70058 153978
rect 75250 148294 75306 148350
rect 75374 148294 75430 148350
rect 75498 148294 75554 148350
rect 75622 148294 75678 148350
rect 75250 148170 75306 148226
rect 75374 148170 75430 148226
rect 75498 148170 75554 148226
rect 75622 148170 75678 148226
rect 75250 148046 75306 148102
rect 75374 148046 75430 148102
rect 75498 148046 75554 148102
rect 75622 148046 75678 148102
rect 75250 147922 75306 147978
rect 75374 147922 75430 147978
rect 75498 147922 75554 147978
rect 75622 147922 75678 147978
rect 60970 136294 61026 136350
rect 61094 136294 61150 136350
rect 61218 136294 61274 136350
rect 61342 136294 61398 136350
rect 60970 136170 61026 136226
rect 61094 136170 61150 136226
rect 61218 136170 61274 136226
rect 61342 136170 61398 136226
rect 60970 136046 61026 136102
rect 61094 136046 61150 136102
rect 61218 136046 61274 136102
rect 61342 136046 61398 136102
rect 60970 135922 61026 135978
rect 61094 135922 61150 135978
rect 61218 135922 61274 135978
rect 61342 135922 61398 135978
rect 69878 136294 69934 136350
rect 70002 136294 70058 136350
rect 69878 136170 69934 136226
rect 70002 136170 70058 136226
rect 69878 136046 69934 136102
rect 70002 136046 70058 136102
rect 69878 135922 69934 135978
rect 70002 135922 70058 135978
rect 75250 130294 75306 130350
rect 75374 130294 75430 130350
rect 75498 130294 75554 130350
rect 75622 130294 75678 130350
rect 75250 130170 75306 130226
rect 75374 130170 75430 130226
rect 75498 130170 75554 130226
rect 75622 130170 75678 130226
rect 75250 130046 75306 130102
rect 75374 130046 75430 130102
rect 75498 130046 75554 130102
rect 75622 130046 75678 130102
rect 75250 129922 75306 129978
rect 75374 129922 75430 129978
rect 75498 129922 75554 129978
rect 75622 129922 75678 129978
rect 60970 118294 61026 118350
rect 61094 118294 61150 118350
rect 61218 118294 61274 118350
rect 61342 118294 61398 118350
rect 60970 118170 61026 118226
rect 61094 118170 61150 118226
rect 61218 118170 61274 118226
rect 61342 118170 61398 118226
rect 60970 118046 61026 118102
rect 61094 118046 61150 118102
rect 61218 118046 61274 118102
rect 61342 118046 61398 118102
rect 60970 117922 61026 117978
rect 61094 117922 61150 117978
rect 61218 117922 61274 117978
rect 61342 117922 61398 117978
rect 69878 118294 69934 118350
rect 70002 118294 70058 118350
rect 69878 118170 69934 118226
rect 70002 118170 70058 118226
rect 69878 118046 69934 118102
rect 70002 118046 70058 118102
rect 69878 117922 69934 117978
rect 70002 117922 70058 117978
rect 75250 112294 75306 112350
rect 75374 112294 75430 112350
rect 75498 112294 75554 112350
rect 75622 112294 75678 112350
rect 75250 112170 75306 112226
rect 75374 112170 75430 112226
rect 75498 112170 75554 112226
rect 75622 112170 75678 112226
rect 75250 112046 75306 112102
rect 75374 112046 75430 112102
rect 75498 112046 75554 112102
rect 75622 112046 75678 112102
rect 75250 111922 75306 111978
rect 75374 111922 75430 111978
rect 75498 111922 75554 111978
rect 75622 111922 75678 111978
rect 60970 100294 61026 100350
rect 61094 100294 61150 100350
rect 61218 100294 61274 100350
rect 61342 100294 61398 100350
rect 60970 100170 61026 100226
rect 61094 100170 61150 100226
rect 61218 100170 61274 100226
rect 61342 100170 61398 100226
rect 60970 100046 61026 100102
rect 61094 100046 61150 100102
rect 61218 100046 61274 100102
rect 61342 100046 61398 100102
rect 60970 99922 61026 99978
rect 61094 99922 61150 99978
rect 61218 99922 61274 99978
rect 61342 99922 61398 99978
rect 69878 100294 69934 100350
rect 70002 100294 70058 100350
rect 69878 100170 69934 100226
rect 70002 100170 70058 100226
rect 69878 100046 69934 100102
rect 70002 100046 70058 100102
rect 69878 99922 69934 99978
rect 70002 99922 70058 99978
rect 75250 94294 75306 94350
rect 75374 94294 75430 94350
rect 75498 94294 75554 94350
rect 75622 94294 75678 94350
rect 75250 94170 75306 94226
rect 75374 94170 75430 94226
rect 75498 94170 75554 94226
rect 75622 94170 75678 94226
rect 75250 94046 75306 94102
rect 75374 94046 75430 94102
rect 75498 94046 75554 94102
rect 75622 94046 75678 94102
rect 75250 93922 75306 93978
rect 75374 93922 75430 93978
rect 75498 93922 75554 93978
rect 75622 93922 75678 93978
rect 60970 82294 61026 82350
rect 61094 82294 61150 82350
rect 61218 82294 61274 82350
rect 61342 82294 61398 82350
rect 60970 82170 61026 82226
rect 61094 82170 61150 82226
rect 61218 82170 61274 82226
rect 61342 82170 61398 82226
rect 60970 82046 61026 82102
rect 61094 82046 61150 82102
rect 61218 82046 61274 82102
rect 61342 82046 61398 82102
rect 60970 81922 61026 81978
rect 61094 81922 61150 81978
rect 61218 81922 61274 81978
rect 61342 81922 61398 81978
rect 69878 82294 69934 82350
rect 70002 82294 70058 82350
rect 69878 82170 69934 82226
rect 70002 82170 70058 82226
rect 69878 82046 69934 82102
rect 70002 82046 70058 82102
rect 69878 81922 69934 81978
rect 70002 81922 70058 81978
rect 75250 76294 75306 76350
rect 75374 76294 75430 76350
rect 75498 76294 75554 76350
rect 75622 76294 75678 76350
rect 75250 76170 75306 76226
rect 75374 76170 75430 76226
rect 75498 76170 75554 76226
rect 75622 76170 75678 76226
rect 75250 76046 75306 76102
rect 75374 76046 75430 76102
rect 75498 76046 75554 76102
rect 75622 76046 75678 76102
rect 75250 75922 75306 75978
rect 75374 75922 75430 75978
rect 75498 75922 75554 75978
rect 75622 75922 75678 75978
rect 60970 64294 61026 64350
rect 61094 64294 61150 64350
rect 61218 64294 61274 64350
rect 61342 64294 61398 64350
rect 60970 64170 61026 64226
rect 61094 64170 61150 64226
rect 61218 64170 61274 64226
rect 61342 64170 61398 64226
rect 60970 64046 61026 64102
rect 61094 64046 61150 64102
rect 61218 64046 61274 64102
rect 61342 64046 61398 64102
rect 60970 63922 61026 63978
rect 61094 63922 61150 63978
rect 61218 63922 61274 63978
rect 61342 63922 61398 63978
rect 69878 64294 69934 64350
rect 70002 64294 70058 64350
rect 69878 64170 69934 64226
rect 70002 64170 70058 64226
rect 69878 64046 69934 64102
rect 70002 64046 70058 64102
rect 69878 63922 69934 63978
rect 70002 63922 70058 63978
rect 75250 58294 75306 58350
rect 75374 58294 75430 58350
rect 75498 58294 75554 58350
rect 75622 58294 75678 58350
rect 75250 58170 75306 58226
rect 75374 58170 75430 58226
rect 75498 58170 75554 58226
rect 75622 58170 75678 58226
rect 75250 58046 75306 58102
rect 75374 58046 75430 58102
rect 75498 58046 75554 58102
rect 75622 58046 75678 58102
rect 75250 57922 75306 57978
rect 75374 57922 75430 57978
rect 75498 57922 75554 57978
rect 75622 57922 75678 57978
rect 60970 46294 61026 46350
rect 61094 46294 61150 46350
rect 61218 46294 61274 46350
rect 61342 46294 61398 46350
rect 60970 46170 61026 46226
rect 61094 46170 61150 46226
rect 61218 46170 61274 46226
rect 61342 46170 61398 46226
rect 60970 46046 61026 46102
rect 61094 46046 61150 46102
rect 61218 46046 61274 46102
rect 61342 46046 61398 46102
rect 60970 45922 61026 45978
rect 61094 45922 61150 45978
rect 61218 45922 61274 45978
rect 61342 45922 61398 45978
rect 69878 46294 69934 46350
rect 70002 46294 70058 46350
rect 69878 46170 69934 46226
rect 70002 46170 70058 46226
rect 69878 46046 69934 46102
rect 70002 46046 70058 46102
rect 69878 45922 69934 45978
rect 70002 45922 70058 45978
rect 60970 28294 61026 28350
rect 61094 28294 61150 28350
rect 61218 28294 61274 28350
rect 61342 28294 61398 28350
rect 60970 28170 61026 28226
rect 61094 28170 61150 28226
rect 61218 28170 61274 28226
rect 61342 28170 61398 28226
rect 60970 28046 61026 28102
rect 61094 28046 61150 28102
rect 61218 28046 61274 28102
rect 61342 28046 61398 28102
rect 60970 27922 61026 27978
rect 61094 27922 61150 27978
rect 61218 27922 61274 27978
rect 61342 27922 61398 27978
rect 60970 10294 61026 10350
rect 61094 10294 61150 10350
rect 61218 10294 61274 10350
rect 61342 10294 61398 10350
rect 60970 10170 61026 10226
rect 61094 10170 61150 10226
rect 61218 10170 61274 10226
rect 61342 10170 61398 10226
rect 60970 10046 61026 10102
rect 61094 10046 61150 10102
rect 61218 10046 61274 10102
rect 61342 10046 61398 10102
rect 60970 9922 61026 9978
rect 61094 9922 61150 9978
rect 61218 9922 61274 9978
rect 61342 9922 61398 9978
rect 60970 -1176 61026 -1120
rect 61094 -1176 61150 -1120
rect 61218 -1176 61274 -1120
rect 61342 -1176 61398 -1120
rect 60970 -1300 61026 -1244
rect 61094 -1300 61150 -1244
rect 61218 -1300 61274 -1244
rect 61342 -1300 61398 -1244
rect 60970 -1424 61026 -1368
rect 61094 -1424 61150 -1368
rect 61218 -1424 61274 -1368
rect 61342 -1424 61398 -1368
rect 60970 -1548 61026 -1492
rect 61094 -1548 61150 -1492
rect 61218 -1548 61274 -1492
rect 61342 -1548 61398 -1492
rect 75250 40294 75306 40350
rect 75374 40294 75430 40350
rect 75498 40294 75554 40350
rect 75622 40294 75678 40350
rect 75250 40170 75306 40226
rect 75374 40170 75430 40226
rect 75498 40170 75554 40226
rect 75622 40170 75678 40226
rect 75250 40046 75306 40102
rect 75374 40046 75430 40102
rect 75498 40046 75554 40102
rect 75622 40046 75678 40102
rect 75250 39922 75306 39978
rect 75374 39922 75430 39978
rect 75498 39922 75554 39978
rect 75622 39922 75678 39978
rect 75250 22294 75306 22350
rect 75374 22294 75430 22350
rect 75498 22294 75554 22350
rect 75622 22294 75678 22350
rect 75250 22170 75306 22226
rect 75374 22170 75430 22226
rect 75498 22170 75554 22226
rect 75622 22170 75678 22226
rect 75250 22046 75306 22102
rect 75374 22046 75430 22102
rect 75498 22046 75554 22102
rect 75622 22046 75678 22102
rect 75250 21922 75306 21978
rect 75374 21922 75430 21978
rect 75498 21922 75554 21978
rect 75622 21922 75678 21978
rect 75250 4294 75306 4350
rect 75374 4294 75430 4350
rect 75498 4294 75554 4350
rect 75622 4294 75678 4350
rect 75250 4170 75306 4226
rect 75374 4170 75430 4226
rect 75498 4170 75554 4226
rect 75622 4170 75678 4226
rect 75250 4046 75306 4102
rect 75374 4046 75430 4102
rect 75498 4046 75554 4102
rect 75622 4046 75678 4102
rect 75250 3922 75306 3978
rect 75374 3922 75430 3978
rect 75498 3922 75554 3978
rect 75622 3922 75678 3978
rect 75250 -216 75306 -160
rect 75374 -216 75430 -160
rect 75498 -216 75554 -160
rect 75622 -216 75678 -160
rect 75250 -340 75306 -284
rect 75374 -340 75430 -284
rect 75498 -340 75554 -284
rect 75622 -340 75678 -284
rect 75250 -464 75306 -408
rect 75374 -464 75430 -408
rect 75498 -464 75554 -408
rect 75622 -464 75678 -408
rect 75250 -588 75306 -532
rect 75374 -588 75430 -532
rect 75498 -588 75554 -532
rect 75622 -588 75678 -532
rect 78970 598116 79026 598172
rect 79094 598116 79150 598172
rect 79218 598116 79274 598172
rect 79342 598116 79398 598172
rect 78970 597992 79026 598048
rect 79094 597992 79150 598048
rect 79218 597992 79274 598048
rect 79342 597992 79398 598048
rect 78970 597868 79026 597924
rect 79094 597868 79150 597924
rect 79218 597868 79274 597924
rect 79342 597868 79398 597924
rect 78970 597744 79026 597800
rect 79094 597744 79150 597800
rect 79218 597744 79274 597800
rect 79342 597744 79398 597800
rect 78970 586294 79026 586350
rect 79094 586294 79150 586350
rect 79218 586294 79274 586350
rect 79342 586294 79398 586350
rect 78970 586170 79026 586226
rect 79094 586170 79150 586226
rect 79218 586170 79274 586226
rect 79342 586170 79398 586226
rect 78970 586046 79026 586102
rect 79094 586046 79150 586102
rect 79218 586046 79274 586102
rect 79342 586046 79398 586102
rect 78970 585922 79026 585978
rect 79094 585922 79150 585978
rect 79218 585922 79274 585978
rect 79342 585922 79398 585978
rect 78970 568294 79026 568350
rect 79094 568294 79150 568350
rect 79218 568294 79274 568350
rect 79342 568294 79398 568350
rect 78970 568170 79026 568226
rect 79094 568170 79150 568226
rect 79218 568170 79274 568226
rect 79342 568170 79398 568226
rect 78970 568046 79026 568102
rect 79094 568046 79150 568102
rect 79218 568046 79274 568102
rect 79342 568046 79398 568102
rect 78970 567922 79026 567978
rect 79094 567922 79150 567978
rect 79218 567922 79274 567978
rect 79342 567922 79398 567978
rect 78970 550294 79026 550350
rect 79094 550294 79150 550350
rect 79218 550294 79274 550350
rect 79342 550294 79398 550350
rect 78970 550170 79026 550226
rect 79094 550170 79150 550226
rect 79218 550170 79274 550226
rect 79342 550170 79398 550226
rect 78970 550046 79026 550102
rect 79094 550046 79150 550102
rect 79218 550046 79274 550102
rect 79342 550046 79398 550102
rect 78970 549922 79026 549978
rect 79094 549922 79150 549978
rect 79218 549922 79274 549978
rect 79342 549922 79398 549978
rect 78970 532294 79026 532350
rect 79094 532294 79150 532350
rect 79218 532294 79274 532350
rect 79342 532294 79398 532350
rect 78970 532170 79026 532226
rect 79094 532170 79150 532226
rect 79218 532170 79274 532226
rect 79342 532170 79398 532226
rect 78970 532046 79026 532102
rect 79094 532046 79150 532102
rect 79218 532046 79274 532102
rect 79342 532046 79398 532102
rect 78970 531922 79026 531978
rect 79094 531922 79150 531978
rect 79218 531922 79274 531978
rect 79342 531922 79398 531978
rect 93250 597156 93306 597212
rect 93374 597156 93430 597212
rect 93498 597156 93554 597212
rect 93622 597156 93678 597212
rect 93250 597032 93306 597088
rect 93374 597032 93430 597088
rect 93498 597032 93554 597088
rect 93622 597032 93678 597088
rect 93250 596908 93306 596964
rect 93374 596908 93430 596964
rect 93498 596908 93554 596964
rect 93622 596908 93678 596964
rect 93250 596784 93306 596840
rect 93374 596784 93430 596840
rect 93498 596784 93554 596840
rect 93622 596784 93678 596840
rect 93250 580294 93306 580350
rect 93374 580294 93430 580350
rect 93498 580294 93554 580350
rect 93622 580294 93678 580350
rect 93250 580170 93306 580226
rect 93374 580170 93430 580226
rect 93498 580170 93554 580226
rect 93622 580170 93678 580226
rect 93250 580046 93306 580102
rect 93374 580046 93430 580102
rect 93498 580046 93554 580102
rect 93622 580046 93678 580102
rect 93250 579922 93306 579978
rect 93374 579922 93430 579978
rect 93498 579922 93554 579978
rect 93622 579922 93678 579978
rect 93250 562294 93306 562350
rect 93374 562294 93430 562350
rect 93498 562294 93554 562350
rect 93622 562294 93678 562350
rect 93250 562170 93306 562226
rect 93374 562170 93430 562226
rect 93498 562170 93554 562226
rect 93622 562170 93678 562226
rect 93250 562046 93306 562102
rect 93374 562046 93430 562102
rect 93498 562046 93554 562102
rect 93622 562046 93678 562102
rect 93250 561922 93306 561978
rect 93374 561922 93430 561978
rect 93498 561922 93554 561978
rect 93622 561922 93678 561978
rect 93250 544294 93306 544350
rect 93374 544294 93430 544350
rect 93498 544294 93554 544350
rect 93622 544294 93678 544350
rect 93250 544170 93306 544226
rect 93374 544170 93430 544226
rect 93498 544170 93554 544226
rect 93622 544170 93678 544226
rect 93250 544046 93306 544102
rect 93374 544046 93430 544102
rect 93498 544046 93554 544102
rect 93622 544046 93678 544102
rect 93250 543922 93306 543978
rect 93374 543922 93430 543978
rect 93498 543922 93554 543978
rect 93622 543922 93678 543978
rect 85238 526237 85294 526293
rect 85362 526237 85418 526293
rect 85238 526113 85294 526169
rect 85362 526113 85418 526169
rect 85238 525989 85294 526045
rect 85362 525989 85418 526045
rect 85238 525865 85294 525921
rect 85362 525865 85418 525921
rect 93250 526294 93306 526350
rect 93374 526294 93430 526350
rect 93498 526294 93554 526350
rect 93622 526294 93678 526350
rect 93250 526170 93306 526226
rect 93374 526170 93430 526226
rect 93498 526170 93554 526226
rect 93622 526170 93678 526226
rect 93250 526046 93306 526102
rect 93374 526046 93430 526102
rect 93498 526046 93554 526102
rect 93622 526046 93678 526102
rect 93250 525922 93306 525978
rect 93374 525922 93430 525978
rect 93498 525922 93554 525978
rect 93622 525922 93678 525978
rect 78970 514294 79026 514350
rect 79094 514294 79150 514350
rect 79218 514294 79274 514350
rect 79342 514294 79398 514350
rect 78970 514170 79026 514226
rect 79094 514170 79150 514226
rect 79218 514170 79274 514226
rect 79342 514170 79398 514226
rect 78970 514046 79026 514102
rect 79094 514046 79150 514102
rect 79218 514046 79274 514102
rect 79342 514046 79398 514102
rect 78970 513922 79026 513978
rect 79094 513922 79150 513978
rect 79218 513922 79274 513978
rect 79342 513922 79398 513978
rect 85238 508294 85294 508350
rect 85362 508294 85418 508350
rect 85238 508170 85294 508226
rect 85362 508170 85418 508226
rect 85238 508046 85294 508102
rect 85362 508046 85418 508102
rect 85238 507922 85294 507978
rect 85362 507922 85418 507978
rect 93250 508294 93306 508350
rect 93374 508294 93430 508350
rect 93498 508294 93554 508350
rect 93622 508294 93678 508350
rect 93250 508170 93306 508226
rect 93374 508170 93430 508226
rect 93498 508170 93554 508226
rect 93622 508170 93678 508226
rect 93250 508046 93306 508102
rect 93374 508046 93430 508102
rect 93498 508046 93554 508102
rect 93622 508046 93678 508102
rect 93250 507922 93306 507978
rect 93374 507922 93430 507978
rect 93498 507922 93554 507978
rect 93622 507922 93678 507978
rect 78970 496294 79026 496350
rect 79094 496294 79150 496350
rect 79218 496294 79274 496350
rect 79342 496294 79398 496350
rect 78970 496170 79026 496226
rect 79094 496170 79150 496226
rect 79218 496170 79274 496226
rect 79342 496170 79398 496226
rect 78970 496046 79026 496102
rect 79094 496046 79150 496102
rect 79218 496046 79274 496102
rect 79342 496046 79398 496102
rect 78970 495922 79026 495978
rect 79094 495922 79150 495978
rect 79218 495922 79274 495978
rect 79342 495922 79398 495978
rect 85238 490294 85294 490350
rect 85362 490294 85418 490350
rect 85238 490170 85294 490226
rect 85362 490170 85418 490226
rect 85238 490046 85294 490102
rect 85362 490046 85418 490102
rect 85238 489922 85294 489978
rect 85362 489922 85418 489978
rect 93250 490294 93306 490350
rect 93374 490294 93430 490350
rect 93498 490294 93554 490350
rect 93622 490294 93678 490350
rect 93250 490170 93306 490226
rect 93374 490170 93430 490226
rect 93498 490170 93554 490226
rect 93622 490170 93678 490226
rect 93250 490046 93306 490102
rect 93374 490046 93430 490102
rect 93498 490046 93554 490102
rect 93622 490046 93678 490102
rect 93250 489922 93306 489978
rect 93374 489922 93430 489978
rect 93498 489922 93554 489978
rect 93622 489922 93678 489978
rect 78970 478294 79026 478350
rect 79094 478294 79150 478350
rect 79218 478294 79274 478350
rect 79342 478294 79398 478350
rect 78970 478170 79026 478226
rect 79094 478170 79150 478226
rect 79218 478170 79274 478226
rect 79342 478170 79398 478226
rect 78970 478046 79026 478102
rect 79094 478046 79150 478102
rect 79218 478046 79274 478102
rect 79342 478046 79398 478102
rect 78970 477922 79026 477978
rect 79094 477922 79150 477978
rect 79218 477922 79274 477978
rect 79342 477922 79398 477978
rect 85238 472294 85294 472350
rect 85362 472294 85418 472350
rect 85238 472170 85294 472226
rect 85362 472170 85418 472226
rect 85238 472046 85294 472102
rect 85362 472046 85418 472102
rect 85238 471922 85294 471978
rect 85362 471922 85418 471978
rect 93250 472294 93306 472350
rect 93374 472294 93430 472350
rect 93498 472294 93554 472350
rect 93622 472294 93678 472350
rect 93250 472170 93306 472226
rect 93374 472170 93430 472226
rect 93498 472170 93554 472226
rect 93622 472170 93678 472226
rect 93250 472046 93306 472102
rect 93374 472046 93430 472102
rect 93498 472046 93554 472102
rect 93622 472046 93678 472102
rect 93250 471922 93306 471978
rect 93374 471922 93430 471978
rect 93498 471922 93554 471978
rect 93622 471922 93678 471978
rect 78970 460294 79026 460350
rect 79094 460294 79150 460350
rect 79218 460294 79274 460350
rect 79342 460294 79398 460350
rect 78970 460170 79026 460226
rect 79094 460170 79150 460226
rect 79218 460170 79274 460226
rect 79342 460170 79398 460226
rect 78970 460046 79026 460102
rect 79094 460046 79150 460102
rect 79218 460046 79274 460102
rect 79342 460046 79398 460102
rect 78970 459922 79026 459978
rect 79094 459922 79150 459978
rect 79218 459922 79274 459978
rect 79342 459922 79398 459978
rect 85238 454294 85294 454350
rect 85362 454294 85418 454350
rect 85238 454170 85294 454226
rect 85362 454170 85418 454226
rect 85238 454046 85294 454102
rect 85362 454046 85418 454102
rect 85238 453922 85294 453978
rect 85362 453922 85418 453978
rect 93250 454294 93306 454350
rect 93374 454294 93430 454350
rect 93498 454294 93554 454350
rect 93622 454294 93678 454350
rect 93250 454170 93306 454226
rect 93374 454170 93430 454226
rect 93498 454170 93554 454226
rect 93622 454170 93678 454226
rect 93250 454046 93306 454102
rect 93374 454046 93430 454102
rect 93498 454046 93554 454102
rect 93622 454046 93678 454102
rect 93250 453922 93306 453978
rect 93374 453922 93430 453978
rect 93498 453922 93554 453978
rect 93622 453922 93678 453978
rect 78970 442294 79026 442350
rect 79094 442294 79150 442350
rect 79218 442294 79274 442350
rect 79342 442294 79398 442350
rect 78970 442170 79026 442226
rect 79094 442170 79150 442226
rect 79218 442170 79274 442226
rect 79342 442170 79398 442226
rect 78970 442046 79026 442102
rect 79094 442046 79150 442102
rect 79218 442046 79274 442102
rect 79342 442046 79398 442102
rect 78970 441922 79026 441978
rect 79094 441922 79150 441978
rect 79218 441922 79274 441978
rect 79342 441922 79398 441978
rect 85238 436294 85294 436350
rect 85362 436294 85418 436350
rect 85238 436170 85294 436226
rect 85362 436170 85418 436226
rect 85238 436046 85294 436102
rect 85362 436046 85418 436102
rect 85238 435922 85294 435978
rect 85362 435922 85418 435978
rect 93250 436294 93306 436350
rect 93374 436294 93430 436350
rect 93498 436294 93554 436350
rect 93622 436294 93678 436350
rect 93250 436170 93306 436226
rect 93374 436170 93430 436226
rect 93498 436170 93554 436226
rect 93622 436170 93678 436226
rect 93250 436046 93306 436102
rect 93374 436046 93430 436102
rect 93498 436046 93554 436102
rect 93622 436046 93678 436102
rect 93250 435922 93306 435978
rect 93374 435922 93430 435978
rect 93498 435922 93554 435978
rect 93622 435922 93678 435978
rect 78970 424294 79026 424350
rect 79094 424294 79150 424350
rect 79218 424294 79274 424350
rect 79342 424294 79398 424350
rect 78970 424170 79026 424226
rect 79094 424170 79150 424226
rect 79218 424170 79274 424226
rect 79342 424170 79398 424226
rect 78970 424046 79026 424102
rect 79094 424046 79150 424102
rect 79218 424046 79274 424102
rect 79342 424046 79398 424102
rect 78970 423922 79026 423978
rect 79094 423922 79150 423978
rect 79218 423922 79274 423978
rect 79342 423922 79398 423978
rect 85238 418294 85294 418350
rect 85362 418294 85418 418350
rect 85238 418170 85294 418226
rect 85362 418170 85418 418226
rect 85238 418046 85294 418102
rect 85362 418046 85418 418102
rect 85238 417922 85294 417978
rect 85362 417922 85418 417978
rect 93250 418294 93306 418350
rect 93374 418294 93430 418350
rect 93498 418294 93554 418350
rect 93622 418294 93678 418350
rect 93250 418170 93306 418226
rect 93374 418170 93430 418226
rect 93498 418170 93554 418226
rect 93622 418170 93678 418226
rect 93250 418046 93306 418102
rect 93374 418046 93430 418102
rect 93498 418046 93554 418102
rect 93622 418046 93678 418102
rect 93250 417922 93306 417978
rect 93374 417922 93430 417978
rect 93498 417922 93554 417978
rect 93622 417922 93678 417978
rect 78970 406294 79026 406350
rect 79094 406294 79150 406350
rect 79218 406294 79274 406350
rect 79342 406294 79398 406350
rect 78970 406170 79026 406226
rect 79094 406170 79150 406226
rect 79218 406170 79274 406226
rect 79342 406170 79398 406226
rect 78970 406046 79026 406102
rect 79094 406046 79150 406102
rect 79218 406046 79274 406102
rect 79342 406046 79398 406102
rect 78970 405922 79026 405978
rect 79094 405922 79150 405978
rect 79218 405922 79274 405978
rect 79342 405922 79398 405978
rect 85238 400294 85294 400350
rect 85362 400294 85418 400350
rect 85238 400170 85294 400226
rect 85362 400170 85418 400226
rect 85238 400046 85294 400102
rect 85362 400046 85418 400102
rect 85238 399922 85294 399978
rect 85362 399922 85418 399978
rect 93250 400294 93306 400350
rect 93374 400294 93430 400350
rect 93498 400294 93554 400350
rect 93622 400294 93678 400350
rect 93250 400170 93306 400226
rect 93374 400170 93430 400226
rect 93498 400170 93554 400226
rect 93622 400170 93678 400226
rect 93250 400046 93306 400102
rect 93374 400046 93430 400102
rect 93498 400046 93554 400102
rect 93622 400046 93678 400102
rect 93250 399922 93306 399978
rect 93374 399922 93430 399978
rect 93498 399922 93554 399978
rect 93622 399922 93678 399978
rect 78970 388294 79026 388350
rect 79094 388294 79150 388350
rect 79218 388294 79274 388350
rect 79342 388294 79398 388350
rect 78970 388170 79026 388226
rect 79094 388170 79150 388226
rect 79218 388170 79274 388226
rect 79342 388170 79398 388226
rect 78970 388046 79026 388102
rect 79094 388046 79150 388102
rect 79218 388046 79274 388102
rect 79342 388046 79398 388102
rect 78970 387922 79026 387978
rect 79094 387922 79150 387978
rect 79218 387922 79274 387978
rect 79342 387922 79398 387978
rect 85238 382294 85294 382350
rect 85362 382294 85418 382350
rect 85238 382170 85294 382226
rect 85362 382170 85418 382226
rect 85238 382046 85294 382102
rect 85362 382046 85418 382102
rect 85238 381922 85294 381978
rect 85362 381922 85418 381978
rect 93250 382294 93306 382350
rect 93374 382294 93430 382350
rect 93498 382294 93554 382350
rect 93622 382294 93678 382350
rect 93250 382170 93306 382226
rect 93374 382170 93430 382226
rect 93498 382170 93554 382226
rect 93622 382170 93678 382226
rect 93250 382046 93306 382102
rect 93374 382046 93430 382102
rect 93498 382046 93554 382102
rect 93622 382046 93678 382102
rect 93250 381922 93306 381978
rect 93374 381922 93430 381978
rect 93498 381922 93554 381978
rect 93622 381922 93678 381978
rect 78970 370294 79026 370350
rect 79094 370294 79150 370350
rect 79218 370294 79274 370350
rect 79342 370294 79398 370350
rect 78970 370170 79026 370226
rect 79094 370170 79150 370226
rect 79218 370170 79274 370226
rect 79342 370170 79398 370226
rect 78970 370046 79026 370102
rect 79094 370046 79150 370102
rect 79218 370046 79274 370102
rect 79342 370046 79398 370102
rect 78970 369922 79026 369978
rect 79094 369922 79150 369978
rect 79218 369922 79274 369978
rect 79342 369922 79398 369978
rect 85238 364294 85294 364350
rect 85362 364294 85418 364350
rect 85238 364170 85294 364226
rect 85362 364170 85418 364226
rect 85238 364046 85294 364102
rect 85362 364046 85418 364102
rect 85238 363922 85294 363978
rect 85362 363922 85418 363978
rect 93250 364294 93306 364350
rect 93374 364294 93430 364350
rect 93498 364294 93554 364350
rect 93622 364294 93678 364350
rect 93250 364170 93306 364226
rect 93374 364170 93430 364226
rect 93498 364170 93554 364226
rect 93622 364170 93678 364226
rect 93250 364046 93306 364102
rect 93374 364046 93430 364102
rect 93498 364046 93554 364102
rect 93622 364046 93678 364102
rect 93250 363922 93306 363978
rect 93374 363922 93430 363978
rect 93498 363922 93554 363978
rect 93622 363922 93678 363978
rect 78970 352294 79026 352350
rect 79094 352294 79150 352350
rect 79218 352294 79274 352350
rect 79342 352294 79398 352350
rect 78970 352170 79026 352226
rect 79094 352170 79150 352226
rect 79218 352170 79274 352226
rect 79342 352170 79398 352226
rect 78970 352046 79026 352102
rect 79094 352046 79150 352102
rect 79218 352046 79274 352102
rect 79342 352046 79398 352102
rect 78970 351922 79026 351978
rect 79094 351922 79150 351978
rect 79218 351922 79274 351978
rect 79342 351922 79398 351978
rect 85238 346294 85294 346350
rect 85362 346294 85418 346350
rect 85238 346170 85294 346226
rect 85362 346170 85418 346226
rect 85238 346046 85294 346102
rect 85362 346046 85418 346102
rect 85238 345922 85294 345978
rect 85362 345922 85418 345978
rect 93250 346294 93306 346350
rect 93374 346294 93430 346350
rect 93498 346294 93554 346350
rect 93622 346294 93678 346350
rect 93250 346170 93306 346226
rect 93374 346170 93430 346226
rect 93498 346170 93554 346226
rect 93622 346170 93678 346226
rect 93250 346046 93306 346102
rect 93374 346046 93430 346102
rect 93498 346046 93554 346102
rect 93622 346046 93678 346102
rect 93250 345922 93306 345978
rect 93374 345922 93430 345978
rect 93498 345922 93554 345978
rect 93622 345922 93678 345978
rect 78970 334294 79026 334350
rect 79094 334294 79150 334350
rect 79218 334294 79274 334350
rect 79342 334294 79398 334350
rect 78970 334170 79026 334226
rect 79094 334170 79150 334226
rect 79218 334170 79274 334226
rect 79342 334170 79398 334226
rect 78970 334046 79026 334102
rect 79094 334046 79150 334102
rect 79218 334046 79274 334102
rect 79342 334046 79398 334102
rect 78970 333922 79026 333978
rect 79094 333922 79150 333978
rect 79218 333922 79274 333978
rect 79342 333922 79398 333978
rect 85238 328294 85294 328350
rect 85362 328294 85418 328350
rect 85238 328170 85294 328226
rect 85362 328170 85418 328226
rect 85238 328046 85294 328102
rect 85362 328046 85418 328102
rect 85238 327922 85294 327978
rect 85362 327922 85418 327978
rect 93250 328294 93306 328350
rect 93374 328294 93430 328350
rect 93498 328294 93554 328350
rect 93622 328294 93678 328350
rect 93250 328170 93306 328226
rect 93374 328170 93430 328226
rect 93498 328170 93554 328226
rect 93622 328170 93678 328226
rect 93250 328046 93306 328102
rect 93374 328046 93430 328102
rect 93498 328046 93554 328102
rect 93622 328046 93678 328102
rect 93250 327922 93306 327978
rect 93374 327922 93430 327978
rect 93498 327922 93554 327978
rect 93622 327922 93678 327978
rect 78970 316294 79026 316350
rect 79094 316294 79150 316350
rect 79218 316294 79274 316350
rect 79342 316294 79398 316350
rect 78970 316170 79026 316226
rect 79094 316170 79150 316226
rect 79218 316170 79274 316226
rect 79342 316170 79398 316226
rect 78970 316046 79026 316102
rect 79094 316046 79150 316102
rect 79218 316046 79274 316102
rect 79342 316046 79398 316102
rect 78970 315922 79026 315978
rect 79094 315922 79150 315978
rect 79218 315922 79274 315978
rect 79342 315922 79398 315978
rect 85238 310294 85294 310350
rect 85362 310294 85418 310350
rect 85238 310170 85294 310226
rect 85362 310170 85418 310226
rect 85238 310046 85294 310102
rect 85362 310046 85418 310102
rect 85238 309922 85294 309978
rect 85362 309922 85418 309978
rect 93250 310294 93306 310350
rect 93374 310294 93430 310350
rect 93498 310294 93554 310350
rect 93622 310294 93678 310350
rect 93250 310170 93306 310226
rect 93374 310170 93430 310226
rect 93498 310170 93554 310226
rect 93622 310170 93678 310226
rect 93250 310046 93306 310102
rect 93374 310046 93430 310102
rect 93498 310046 93554 310102
rect 93622 310046 93678 310102
rect 93250 309922 93306 309978
rect 93374 309922 93430 309978
rect 93498 309922 93554 309978
rect 93622 309922 93678 309978
rect 78970 298294 79026 298350
rect 79094 298294 79150 298350
rect 79218 298294 79274 298350
rect 79342 298294 79398 298350
rect 78970 298170 79026 298226
rect 79094 298170 79150 298226
rect 79218 298170 79274 298226
rect 79342 298170 79398 298226
rect 78970 298046 79026 298102
rect 79094 298046 79150 298102
rect 79218 298046 79274 298102
rect 79342 298046 79398 298102
rect 78970 297922 79026 297978
rect 79094 297922 79150 297978
rect 79218 297922 79274 297978
rect 79342 297922 79398 297978
rect 85238 292294 85294 292350
rect 85362 292294 85418 292350
rect 85238 292170 85294 292226
rect 85362 292170 85418 292226
rect 85238 292046 85294 292102
rect 85362 292046 85418 292102
rect 85238 291922 85294 291978
rect 85362 291922 85418 291978
rect 93250 292294 93306 292350
rect 93374 292294 93430 292350
rect 93498 292294 93554 292350
rect 93622 292294 93678 292350
rect 93250 292170 93306 292226
rect 93374 292170 93430 292226
rect 93498 292170 93554 292226
rect 93622 292170 93678 292226
rect 93250 292046 93306 292102
rect 93374 292046 93430 292102
rect 93498 292046 93554 292102
rect 93622 292046 93678 292102
rect 93250 291922 93306 291978
rect 93374 291922 93430 291978
rect 93498 291922 93554 291978
rect 93622 291922 93678 291978
rect 78970 280294 79026 280350
rect 79094 280294 79150 280350
rect 79218 280294 79274 280350
rect 79342 280294 79398 280350
rect 78970 280170 79026 280226
rect 79094 280170 79150 280226
rect 79218 280170 79274 280226
rect 79342 280170 79398 280226
rect 78970 280046 79026 280102
rect 79094 280046 79150 280102
rect 79218 280046 79274 280102
rect 79342 280046 79398 280102
rect 78970 279922 79026 279978
rect 79094 279922 79150 279978
rect 79218 279922 79274 279978
rect 79342 279922 79398 279978
rect 85238 274294 85294 274350
rect 85362 274294 85418 274350
rect 85238 274170 85294 274226
rect 85362 274170 85418 274226
rect 85238 274046 85294 274102
rect 85362 274046 85418 274102
rect 85238 273922 85294 273978
rect 85362 273922 85418 273978
rect 93250 274294 93306 274350
rect 93374 274294 93430 274350
rect 93498 274294 93554 274350
rect 93622 274294 93678 274350
rect 93250 274170 93306 274226
rect 93374 274170 93430 274226
rect 93498 274170 93554 274226
rect 93622 274170 93678 274226
rect 93250 274046 93306 274102
rect 93374 274046 93430 274102
rect 93498 274046 93554 274102
rect 93622 274046 93678 274102
rect 93250 273922 93306 273978
rect 93374 273922 93430 273978
rect 93498 273922 93554 273978
rect 93622 273922 93678 273978
rect 78970 262294 79026 262350
rect 79094 262294 79150 262350
rect 79218 262294 79274 262350
rect 79342 262294 79398 262350
rect 78970 262170 79026 262226
rect 79094 262170 79150 262226
rect 79218 262170 79274 262226
rect 79342 262170 79398 262226
rect 78970 262046 79026 262102
rect 79094 262046 79150 262102
rect 79218 262046 79274 262102
rect 79342 262046 79398 262102
rect 78970 261922 79026 261978
rect 79094 261922 79150 261978
rect 79218 261922 79274 261978
rect 79342 261922 79398 261978
rect 85238 256294 85294 256350
rect 85362 256294 85418 256350
rect 85238 256170 85294 256226
rect 85362 256170 85418 256226
rect 85238 256046 85294 256102
rect 85362 256046 85418 256102
rect 85238 255922 85294 255978
rect 85362 255922 85418 255978
rect 93250 256294 93306 256350
rect 93374 256294 93430 256350
rect 93498 256294 93554 256350
rect 93622 256294 93678 256350
rect 93250 256170 93306 256226
rect 93374 256170 93430 256226
rect 93498 256170 93554 256226
rect 93622 256170 93678 256226
rect 93250 256046 93306 256102
rect 93374 256046 93430 256102
rect 93498 256046 93554 256102
rect 93622 256046 93678 256102
rect 93250 255922 93306 255978
rect 93374 255922 93430 255978
rect 93498 255922 93554 255978
rect 93622 255922 93678 255978
rect 78970 244294 79026 244350
rect 79094 244294 79150 244350
rect 79218 244294 79274 244350
rect 79342 244294 79398 244350
rect 78970 244170 79026 244226
rect 79094 244170 79150 244226
rect 79218 244170 79274 244226
rect 79342 244170 79398 244226
rect 78970 244046 79026 244102
rect 79094 244046 79150 244102
rect 79218 244046 79274 244102
rect 79342 244046 79398 244102
rect 78970 243922 79026 243978
rect 79094 243922 79150 243978
rect 79218 243922 79274 243978
rect 79342 243922 79398 243978
rect 85238 238294 85294 238350
rect 85362 238294 85418 238350
rect 85238 238170 85294 238226
rect 85362 238170 85418 238226
rect 85238 238046 85294 238102
rect 85362 238046 85418 238102
rect 85238 237922 85294 237978
rect 85362 237922 85418 237978
rect 93250 238294 93306 238350
rect 93374 238294 93430 238350
rect 93498 238294 93554 238350
rect 93622 238294 93678 238350
rect 93250 238170 93306 238226
rect 93374 238170 93430 238226
rect 93498 238170 93554 238226
rect 93622 238170 93678 238226
rect 93250 238046 93306 238102
rect 93374 238046 93430 238102
rect 93498 238046 93554 238102
rect 93622 238046 93678 238102
rect 93250 237922 93306 237978
rect 93374 237922 93430 237978
rect 93498 237922 93554 237978
rect 93622 237922 93678 237978
rect 78970 226294 79026 226350
rect 79094 226294 79150 226350
rect 79218 226294 79274 226350
rect 79342 226294 79398 226350
rect 78970 226170 79026 226226
rect 79094 226170 79150 226226
rect 79218 226170 79274 226226
rect 79342 226170 79398 226226
rect 78970 226046 79026 226102
rect 79094 226046 79150 226102
rect 79218 226046 79274 226102
rect 79342 226046 79398 226102
rect 78970 225922 79026 225978
rect 79094 225922 79150 225978
rect 79218 225922 79274 225978
rect 79342 225922 79398 225978
rect 85238 220294 85294 220350
rect 85362 220294 85418 220350
rect 85238 220170 85294 220226
rect 85362 220170 85418 220226
rect 85238 220046 85294 220102
rect 85362 220046 85418 220102
rect 85238 219922 85294 219978
rect 85362 219922 85418 219978
rect 93250 220294 93306 220350
rect 93374 220294 93430 220350
rect 93498 220294 93554 220350
rect 93622 220294 93678 220350
rect 93250 220170 93306 220226
rect 93374 220170 93430 220226
rect 93498 220170 93554 220226
rect 93622 220170 93678 220226
rect 93250 220046 93306 220102
rect 93374 220046 93430 220102
rect 93498 220046 93554 220102
rect 93622 220046 93678 220102
rect 93250 219922 93306 219978
rect 93374 219922 93430 219978
rect 93498 219922 93554 219978
rect 93622 219922 93678 219978
rect 78970 208294 79026 208350
rect 79094 208294 79150 208350
rect 79218 208294 79274 208350
rect 79342 208294 79398 208350
rect 78970 208170 79026 208226
rect 79094 208170 79150 208226
rect 79218 208170 79274 208226
rect 79342 208170 79398 208226
rect 78970 208046 79026 208102
rect 79094 208046 79150 208102
rect 79218 208046 79274 208102
rect 79342 208046 79398 208102
rect 78970 207922 79026 207978
rect 79094 207922 79150 207978
rect 79218 207922 79274 207978
rect 79342 207922 79398 207978
rect 85238 202294 85294 202350
rect 85362 202294 85418 202350
rect 85238 202170 85294 202226
rect 85362 202170 85418 202226
rect 85238 202046 85294 202102
rect 85362 202046 85418 202102
rect 85238 201922 85294 201978
rect 85362 201922 85418 201978
rect 93250 202294 93306 202350
rect 93374 202294 93430 202350
rect 93498 202294 93554 202350
rect 93622 202294 93678 202350
rect 93250 202170 93306 202226
rect 93374 202170 93430 202226
rect 93498 202170 93554 202226
rect 93622 202170 93678 202226
rect 93250 202046 93306 202102
rect 93374 202046 93430 202102
rect 93498 202046 93554 202102
rect 93622 202046 93678 202102
rect 93250 201922 93306 201978
rect 93374 201922 93430 201978
rect 93498 201922 93554 201978
rect 93622 201922 93678 201978
rect 78970 190294 79026 190350
rect 79094 190294 79150 190350
rect 79218 190294 79274 190350
rect 79342 190294 79398 190350
rect 78970 190170 79026 190226
rect 79094 190170 79150 190226
rect 79218 190170 79274 190226
rect 79342 190170 79398 190226
rect 78970 190046 79026 190102
rect 79094 190046 79150 190102
rect 79218 190046 79274 190102
rect 79342 190046 79398 190102
rect 78970 189922 79026 189978
rect 79094 189922 79150 189978
rect 79218 189922 79274 189978
rect 79342 189922 79398 189978
rect 85238 184294 85294 184350
rect 85362 184294 85418 184350
rect 85238 184170 85294 184226
rect 85362 184170 85418 184226
rect 85238 184046 85294 184102
rect 85362 184046 85418 184102
rect 85238 183922 85294 183978
rect 85362 183922 85418 183978
rect 93250 184294 93306 184350
rect 93374 184294 93430 184350
rect 93498 184294 93554 184350
rect 93622 184294 93678 184350
rect 93250 184170 93306 184226
rect 93374 184170 93430 184226
rect 93498 184170 93554 184226
rect 93622 184170 93678 184226
rect 93250 184046 93306 184102
rect 93374 184046 93430 184102
rect 93498 184046 93554 184102
rect 93622 184046 93678 184102
rect 93250 183922 93306 183978
rect 93374 183922 93430 183978
rect 93498 183922 93554 183978
rect 93622 183922 93678 183978
rect 78970 172294 79026 172350
rect 79094 172294 79150 172350
rect 79218 172294 79274 172350
rect 79342 172294 79398 172350
rect 78970 172170 79026 172226
rect 79094 172170 79150 172226
rect 79218 172170 79274 172226
rect 79342 172170 79398 172226
rect 78970 172046 79026 172102
rect 79094 172046 79150 172102
rect 79218 172046 79274 172102
rect 79342 172046 79398 172102
rect 78970 171922 79026 171978
rect 79094 171922 79150 171978
rect 79218 171922 79274 171978
rect 79342 171922 79398 171978
rect 85238 166294 85294 166350
rect 85362 166294 85418 166350
rect 85238 166170 85294 166226
rect 85362 166170 85418 166226
rect 85238 166046 85294 166102
rect 85362 166046 85418 166102
rect 85238 165922 85294 165978
rect 85362 165922 85418 165978
rect 93250 166294 93306 166350
rect 93374 166294 93430 166350
rect 93498 166294 93554 166350
rect 93622 166294 93678 166350
rect 93250 166170 93306 166226
rect 93374 166170 93430 166226
rect 93498 166170 93554 166226
rect 93622 166170 93678 166226
rect 93250 166046 93306 166102
rect 93374 166046 93430 166102
rect 93498 166046 93554 166102
rect 93622 166046 93678 166102
rect 93250 165922 93306 165978
rect 93374 165922 93430 165978
rect 93498 165922 93554 165978
rect 93622 165922 93678 165978
rect 78970 154294 79026 154350
rect 79094 154294 79150 154350
rect 79218 154294 79274 154350
rect 79342 154294 79398 154350
rect 78970 154170 79026 154226
rect 79094 154170 79150 154226
rect 79218 154170 79274 154226
rect 79342 154170 79398 154226
rect 78970 154046 79026 154102
rect 79094 154046 79150 154102
rect 79218 154046 79274 154102
rect 79342 154046 79398 154102
rect 78970 153922 79026 153978
rect 79094 153922 79150 153978
rect 79218 153922 79274 153978
rect 79342 153922 79398 153978
rect 85238 148294 85294 148350
rect 85362 148294 85418 148350
rect 85238 148170 85294 148226
rect 85362 148170 85418 148226
rect 85238 148046 85294 148102
rect 85362 148046 85418 148102
rect 85238 147922 85294 147978
rect 85362 147922 85418 147978
rect 93250 148294 93306 148350
rect 93374 148294 93430 148350
rect 93498 148294 93554 148350
rect 93622 148294 93678 148350
rect 93250 148170 93306 148226
rect 93374 148170 93430 148226
rect 93498 148170 93554 148226
rect 93622 148170 93678 148226
rect 93250 148046 93306 148102
rect 93374 148046 93430 148102
rect 93498 148046 93554 148102
rect 93622 148046 93678 148102
rect 93250 147922 93306 147978
rect 93374 147922 93430 147978
rect 93498 147922 93554 147978
rect 93622 147922 93678 147978
rect 78970 136294 79026 136350
rect 79094 136294 79150 136350
rect 79218 136294 79274 136350
rect 79342 136294 79398 136350
rect 78970 136170 79026 136226
rect 79094 136170 79150 136226
rect 79218 136170 79274 136226
rect 79342 136170 79398 136226
rect 78970 136046 79026 136102
rect 79094 136046 79150 136102
rect 79218 136046 79274 136102
rect 79342 136046 79398 136102
rect 78970 135922 79026 135978
rect 79094 135922 79150 135978
rect 79218 135922 79274 135978
rect 79342 135922 79398 135978
rect 85238 130294 85294 130350
rect 85362 130294 85418 130350
rect 85238 130170 85294 130226
rect 85362 130170 85418 130226
rect 85238 130046 85294 130102
rect 85362 130046 85418 130102
rect 85238 129922 85294 129978
rect 85362 129922 85418 129978
rect 93250 130294 93306 130350
rect 93374 130294 93430 130350
rect 93498 130294 93554 130350
rect 93622 130294 93678 130350
rect 93250 130170 93306 130226
rect 93374 130170 93430 130226
rect 93498 130170 93554 130226
rect 93622 130170 93678 130226
rect 93250 130046 93306 130102
rect 93374 130046 93430 130102
rect 93498 130046 93554 130102
rect 93622 130046 93678 130102
rect 93250 129922 93306 129978
rect 93374 129922 93430 129978
rect 93498 129922 93554 129978
rect 93622 129922 93678 129978
rect 78970 118294 79026 118350
rect 79094 118294 79150 118350
rect 79218 118294 79274 118350
rect 79342 118294 79398 118350
rect 78970 118170 79026 118226
rect 79094 118170 79150 118226
rect 79218 118170 79274 118226
rect 79342 118170 79398 118226
rect 78970 118046 79026 118102
rect 79094 118046 79150 118102
rect 79218 118046 79274 118102
rect 79342 118046 79398 118102
rect 78970 117922 79026 117978
rect 79094 117922 79150 117978
rect 79218 117922 79274 117978
rect 79342 117922 79398 117978
rect 85238 112294 85294 112350
rect 85362 112294 85418 112350
rect 85238 112170 85294 112226
rect 85362 112170 85418 112226
rect 85238 112046 85294 112102
rect 85362 112046 85418 112102
rect 85238 111922 85294 111978
rect 85362 111922 85418 111978
rect 93250 112294 93306 112350
rect 93374 112294 93430 112350
rect 93498 112294 93554 112350
rect 93622 112294 93678 112350
rect 93250 112170 93306 112226
rect 93374 112170 93430 112226
rect 93498 112170 93554 112226
rect 93622 112170 93678 112226
rect 93250 112046 93306 112102
rect 93374 112046 93430 112102
rect 93498 112046 93554 112102
rect 93622 112046 93678 112102
rect 93250 111922 93306 111978
rect 93374 111922 93430 111978
rect 93498 111922 93554 111978
rect 93622 111922 93678 111978
rect 78970 100294 79026 100350
rect 79094 100294 79150 100350
rect 79218 100294 79274 100350
rect 79342 100294 79398 100350
rect 78970 100170 79026 100226
rect 79094 100170 79150 100226
rect 79218 100170 79274 100226
rect 79342 100170 79398 100226
rect 78970 100046 79026 100102
rect 79094 100046 79150 100102
rect 79218 100046 79274 100102
rect 79342 100046 79398 100102
rect 78970 99922 79026 99978
rect 79094 99922 79150 99978
rect 79218 99922 79274 99978
rect 79342 99922 79398 99978
rect 85238 94294 85294 94350
rect 85362 94294 85418 94350
rect 85238 94170 85294 94226
rect 85362 94170 85418 94226
rect 85238 94046 85294 94102
rect 85362 94046 85418 94102
rect 85238 93922 85294 93978
rect 85362 93922 85418 93978
rect 93250 94294 93306 94350
rect 93374 94294 93430 94350
rect 93498 94294 93554 94350
rect 93622 94294 93678 94350
rect 93250 94170 93306 94226
rect 93374 94170 93430 94226
rect 93498 94170 93554 94226
rect 93622 94170 93678 94226
rect 93250 94046 93306 94102
rect 93374 94046 93430 94102
rect 93498 94046 93554 94102
rect 93622 94046 93678 94102
rect 93250 93922 93306 93978
rect 93374 93922 93430 93978
rect 93498 93922 93554 93978
rect 93622 93922 93678 93978
rect 78970 82294 79026 82350
rect 79094 82294 79150 82350
rect 79218 82294 79274 82350
rect 79342 82294 79398 82350
rect 78970 82170 79026 82226
rect 79094 82170 79150 82226
rect 79218 82170 79274 82226
rect 79342 82170 79398 82226
rect 78970 82046 79026 82102
rect 79094 82046 79150 82102
rect 79218 82046 79274 82102
rect 79342 82046 79398 82102
rect 78970 81922 79026 81978
rect 79094 81922 79150 81978
rect 79218 81922 79274 81978
rect 79342 81922 79398 81978
rect 85238 76294 85294 76350
rect 85362 76294 85418 76350
rect 85238 76170 85294 76226
rect 85362 76170 85418 76226
rect 85238 76046 85294 76102
rect 85362 76046 85418 76102
rect 85238 75922 85294 75978
rect 85362 75922 85418 75978
rect 93250 76294 93306 76350
rect 93374 76294 93430 76350
rect 93498 76294 93554 76350
rect 93622 76294 93678 76350
rect 93250 76170 93306 76226
rect 93374 76170 93430 76226
rect 93498 76170 93554 76226
rect 93622 76170 93678 76226
rect 93250 76046 93306 76102
rect 93374 76046 93430 76102
rect 93498 76046 93554 76102
rect 93622 76046 93678 76102
rect 93250 75922 93306 75978
rect 93374 75922 93430 75978
rect 93498 75922 93554 75978
rect 93622 75922 93678 75978
rect 78970 64294 79026 64350
rect 79094 64294 79150 64350
rect 79218 64294 79274 64350
rect 79342 64294 79398 64350
rect 78970 64170 79026 64226
rect 79094 64170 79150 64226
rect 79218 64170 79274 64226
rect 79342 64170 79398 64226
rect 78970 64046 79026 64102
rect 79094 64046 79150 64102
rect 79218 64046 79274 64102
rect 79342 64046 79398 64102
rect 78970 63922 79026 63978
rect 79094 63922 79150 63978
rect 79218 63922 79274 63978
rect 79342 63922 79398 63978
rect 85238 58294 85294 58350
rect 85362 58294 85418 58350
rect 85238 58170 85294 58226
rect 85362 58170 85418 58226
rect 85238 58046 85294 58102
rect 85362 58046 85418 58102
rect 85238 57922 85294 57978
rect 85362 57922 85418 57978
rect 93250 58294 93306 58350
rect 93374 58294 93430 58350
rect 93498 58294 93554 58350
rect 93622 58294 93678 58350
rect 93250 58170 93306 58226
rect 93374 58170 93430 58226
rect 93498 58170 93554 58226
rect 93622 58170 93678 58226
rect 93250 58046 93306 58102
rect 93374 58046 93430 58102
rect 93498 58046 93554 58102
rect 93622 58046 93678 58102
rect 93250 57922 93306 57978
rect 93374 57922 93430 57978
rect 93498 57922 93554 57978
rect 93622 57922 93678 57978
rect 78970 46294 79026 46350
rect 79094 46294 79150 46350
rect 79218 46294 79274 46350
rect 79342 46294 79398 46350
rect 78970 46170 79026 46226
rect 79094 46170 79150 46226
rect 79218 46170 79274 46226
rect 79342 46170 79398 46226
rect 78970 46046 79026 46102
rect 79094 46046 79150 46102
rect 79218 46046 79274 46102
rect 79342 46046 79398 46102
rect 78970 45922 79026 45978
rect 79094 45922 79150 45978
rect 79218 45922 79274 45978
rect 79342 45922 79398 45978
rect 85238 40294 85294 40350
rect 85362 40294 85418 40350
rect 85238 40170 85294 40226
rect 85362 40170 85418 40226
rect 85238 40046 85294 40102
rect 85362 40046 85418 40102
rect 85238 39922 85294 39978
rect 85362 39922 85418 39978
rect 93250 40294 93306 40350
rect 93374 40294 93430 40350
rect 93498 40294 93554 40350
rect 93622 40294 93678 40350
rect 93250 40170 93306 40226
rect 93374 40170 93430 40226
rect 93498 40170 93554 40226
rect 93622 40170 93678 40226
rect 93250 40046 93306 40102
rect 93374 40046 93430 40102
rect 93498 40046 93554 40102
rect 93622 40046 93678 40102
rect 93250 39922 93306 39978
rect 93374 39922 93430 39978
rect 93498 39922 93554 39978
rect 93622 39922 93678 39978
rect 78970 28294 79026 28350
rect 79094 28294 79150 28350
rect 79218 28294 79274 28350
rect 79342 28294 79398 28350
rect 78970 28170 79026 28226
rect 79094 28170 79150 28226
rect 79218 28170 79274 28226
rect 79342 28170 79398 28226
rect 78970 28046 79026 28102
rect 79094 28046 79150 28102
rect 79218 28046 79274 28102
rect 79342 28046 79398 28102
rect 78970 27922 79026 27978
rect 79094 27922 79150 27978
rect 79218 27922 79274 27978
rect 79342 27922 79398 27978
rect 78970 10294 79026 10350
rect 79094 10294 79150 10350
rect 79218 10294 79274 10350
rect 79342 10294 79398 10350
rect 78970 10170 79026 10226
rect 79094 10170 79150 10226
rect 79218 10170 79274 10226
rect 79342 10170 79398 10226
rect 78970 10046 79026 10102
rect 79094 10046 79150 10102
rect 79218 10046 79274 10102
rect 79342 10046 79398 10102
rect 78970 9922 79026 9978
rect 79094 9922 79150 9978
rect 79218 9922 79274 9978
rect 79342 9922 79398 9978
rect 78970 -1176 79026 -1120
rect 79094 -1176 79150 -1120
rect 79218 -1176 79274 -1120
rect 79342 -1176 79398 -1120
rect 78970 -1300 79026 -1244
rect 79094 -1300 79150 -1244
rect 79218 -1300 79274 -1244
rect 79342 -1300 79398 -1244
rect 78970 -1424 79026 -1368
rect 79094 -1424 79150 -1368
rect 79218 -1424 79274 -1368
rect 79342 -1424 79398 -1368
rect 78970 -1548 79026 -1492
rect 79094 -1548 79150 -1492
rect 79218 -1548 79274 -1492
rect 79342 -1548 79398 -1492
rect 93250 22294 93306 22350
rect 93374 22294 93430 22350
rect 93498 22294 93554 22350
rect 93622 22294 93678 22350
rect 93250 22170 93306 22226
rect 93374 22170 93430 22226
rect 93498 22170 93554 22226
rect 93622 22170 93678 22226
rect 93250 22046 93306 22102
rect 93374 22046 93430 22102
rect 93498 22046 93554 22102
rect 93622 22046 93678 22102
rect 93250 21922 93306 21978
rect 93374 21922 93430 21978
rect 93498 21922 93554 21978
rect 93622 21922 93678 21978
rect 93250 4294 93306 4350
rect 93374 4294 93430 4350
rect 93498 4294 93554 4350
rect 93622 4294 93678 4350
rect 93250 4170 93306 4226
rect 93374 4170 93430 4226
rect 93498 4170 93554 4226
rect 93622 4170 93678 4226
rect 93250 4046 93306 4102
rect 93374 4046 93430 4102
rect 93498 4046 93554 4102
rect 93622 4046 93678 4102
rect 93250 3922 93306 3978
rect 93374 3922 93430 3978
rect 93498 3922 93554 3978
rect 93622 3922 93678 3978
rect 93250 -216 93306 -160
rect 93374 -216 93430 -160
rect 93498 -216 93554 -160
rect 93622 -216 93678 -160
rect 93250 -340 93306 -284
rect 93374 -340 93430 -284
rect 93498 -340 93554 -284
rect 93622 -340 93678 -284
rect 93250 -464 93306 -408
rect 93374 -464 93430 -408
rect 93498 -464 93554 -408
rect 93622 -464 93678 -408
rect 93250 -588 93306 -532
rect 93374 -588 93430 -532
rect 93498 -588 93554 -532
rect 93622 -588 93678 -532
rect 96970 598116 97026 598172
rect 97094 598116 97150 598172
rect 97218 598116 97274 598172
rect 97342 598116 97398 598172
rect 96970 597992 97026 598048
rect 97094 597992 97150 598048
rect 97218 597992 97274 598048
rect 97342 597992 97398 598048
rect 96970 597868 97026 597924
rect 97094 597868 97150 597924
rect 97218 597868 97274 597924
rect 97342 597868 97398 597924
rect 96970 597744 97026 597800
rect 97094 597744 97150 597800
rect 97218 597744 97274 597800
rect 97342 597744 97398 597800
rect 96970 586294 97026 586350
rect 97094 586294 97150 586350
rect 97218 586294 97274 586350
rect 97342 586294 97398 586350
rect 96970 586170 97026 586226
rect 97094 586170 97150 586226
rect 97218 586170 97274 586226
rect 97342 586170 97398 586226
rect 96970 586046 97026 586102
rect 97094 586046 97150 586102
rect 97218 586046 97274 586102
rect 97342 586046 97398 586102
rect 96970 585922 97026 585978
rect 97094 585922 97150 585978
rect 97218 585922 97274 585978
rect 97342 585922 97398 585978
rect 96970 568294 97026 568350
rect 97094 568294 97150 568350
rect 97218 568294 97274 568350
rect 97342 568294 97398 568350
rect 96970 568170 97026 568226
rect 97094 568170 97150 568226
rect 97218 568170 97274 568226
rect 97342 568170 97398 568226
rect 96970 568046 97026 568102
rect 97094 568046 97150 568102
rect 97218 568046 97274 568102
rect 97342 568046 97398 568102
rect 96970 567922 97026 567978
rect 97094 567922 97150 567978
rect 97218 567922 97274 567978
rect 97342 567922 97398 567978
rect 96970 550294 97026 550350
rect 97094 550294 97150 550350
rect 97218 550294 97274 550350
rect 97342 550294 97398 550350
rect 96970 550170 97026 550226
rect 97094 550170 97150 550226
rect 97218 550170 97274 550226
rect 97342 550170 97398 550226
rect 96970 550046 97026 550102
rect 97094 550046 97150 550102
rect 97218 550046 97274 550102
rect 97342 550046 97398 550102
rect 96970 549922 97026 549978
rect 97094 549922 97150 549978
rect 97218 549922 97274 549978
rect 97342 549922 97398 549978
rect 96970 532294 97026 532350
rect 97094 532294 97150 532350
rect 97218 532294 97274 532350
rect 97342 532294 97398 532350
rect 96970 532170 97026 532226
rect 97094 532170 97150 532226
rect 97218 532170 97274 532226
rect 97342 532170 97398 532226
rect 96970 532046 97026 532102
rect 97094 532046 97150 532102
rect 97218 532046 97274 532102
rect 97342 532046 97398 532102
rect 96970 531922 97026 531978
rect 97094 531922 97150 531978
rect 97218 531922 97274 531978
rect 97342 531922 97398 531978
rect 111250 597156 111306 597212
rect 111374 597156 111430 597212
rect 111498 597156 111554 597212
rect 111622 597156 111678 597212
rect 111250 597032 111306 597088
rect 111374 597032 111430 597088
rect 111498 597032 111554 597088
rect 111622 597032 111678 597088
rect 111250 596908 111306 596964
rect 111374 596908 111430 596964
rect 111498 596908 111554 596964
rect 111622 596908 111678 596964
rect 111250 596784 111306 596840
rect 111374 596784 111430 596840
rect 111498 596784 111554 596840
rect 111622 596784 111678 596840
rect 111250 580294 111306 580350
rect 111374 580294 111430 580350
rect 111498 580294 111554 580350
rect 111622 580294 111678 580350
rect 111250 580170 111306 580226
rect 111374 580170 111430 580226
rect 111498 580170 111554 580226
rect 111622 580170 111678 580226
rect 111250 580046 111306 580102
rect 111374 580046 111430 580102
rect 111498 580046 111554 580102
rect 111622 580046 111678 580102
rect 111250 579922 111306 579978
rect 111374 579922 111430 579978
rect 111498 579922 111554 579978
rect 111622 579922 111678 579978
rect 111250 562294 111306 562350
rect 111374 562294 111430 562350
rect 111498 562294 111554 562350
rect 111622 562294 111678 562350
rect 111250 562170 111306 562226
rect 111374 562170 111430 562226
rect 111498 562170 111554 562226
rect 111622 562170 111678 562226
rect 111250 562046 111306 562102
rect 111374 562046 111430 562102
rect 111498 562046 111554 562102
rect 111622 562046 111678 562102
rect 111250 561922 111306 561978
rect 111374 561922 111430 561978
rect 111498 561922 111554 561978
rect 111622 561922 111678 561978
rect 111250 544294 111306 544350
rect 111374 544294 111430 544350
rect 111498 544294 111554 544350
rect 111622 544294 111678 544350
rect 111250 544170 111306 544226
rect 111374 544170 111430 544226
rect 111498 544170 111554 544226
rect 111622 544170 111678 544226
rect 111250 544046 111306 544102
rect 111374 544046 111430 544102
rect 111498 544046 111554 544102
rect 111622 544046 111678 544102
rect 111250 543922 111306 543978
rect 111374 543922 111430 543978
rect 111498 543922 111554 543978
rect 111622 543922 111678 543978
rect 114970 598116 115026 598172
rect 115094 598116 115150 598172
rect 115218 598116 115274 598172
rect 115342 598116 115398 598172
rect 114970 597992 115026 598048
rect 115094 597992 115150 598048
rect 115218 597992 115274 598048
rect 115342 597992 115398 598048
rect 114970 597868 115026 597924
rect 115094 597868 115150 597924
rect 115218 597868 115274 597924
rect 115342 597868 115398 597924
rect 114970 597744 115026 597800
rect 115094 597744 115150 597800
rect 115218 597744 115274 597800
rect 115342 597744 115398 597800
rect 114970 586294 115026 586350
rect 115094 586294 115150 586350
rect 115218 586294 115274 586350
rect 115342 586294 115398 586350
rect 114970 586170 115026 586226
rect 115094 586170 115150 586226
rect 115218 586170 115274 586226
rect 115342 586170 115398 586226
rect 114970 586046 115026 586102
rect 115094 586046 115150 586102
rect 115218 586046 115274 586102
rect 115342 586046 115398 586102
rect 114970 585922 115026 585978
rect 115094 585922 115150 585978
rect 115218 585922 115274 585978
rect 115342 585922 115398 585978
rect 114970 568294 115026 568350
rect 115094 568294 115150 568350
rect 115218 568294 115274 568350
rect 115342 568294 115398 568350
rect 114970 568170 115026 568226
rect 115094 568170 115150 568226
rect 115218 568170 115274 568226
rect 115342 568170 115398 568226
rect 114970 568046 115026 568102
rect 115094 568046 115150 568102
rect 115218 568046 115274 568102
rect 115342 568046 115398 568102
rect 114970 567922 115026 567978
rect 115094 567922 115150 567978
rect 115218 567922 115274 567978
rect 115342 567922 115398 567978
rect 114970 550294 115026 550350
rect 115094 550294 115150 550350
rect 115218 550294 115274 550350
rect 115342 550294 115398 550350
rect 114970 550170 115026 550226
rect 115094 550170 115150 550226
rect 115218 550170 115274 550226
rect 115342 550170 115398 550226
rect 114970 550046 115026 550102
rect 115094 550046 115150 550102
rect 115218 550046 115274 550102
rect 115342 550046 115398 550102
rect 114970 549922 115026 549978
rect 115094 549922 115150 549978
rect 115218 549922 115274 549978
rect 115342 549922 115398 549978
rect 114970 532294 115026 532350
rect 115094 532294 115150 532350
rect 115218 532294 115274 532350
rect 115342 532294 115398 532350
rect 114970 532170 115026 532226
rect 115094 532170 115150 532226
rect 115218 532170 115274 532226
rect 115342 532170 115398 532226
rect 114970 532046 115026 532102
rect 115094 532046 115150 532102
rect 115218 532046 115274 532102
rect 115342 532046 115398 532102
rect 114970 531922 115026 531978
rect 115094 531922 115150 531978
rect 115218 531922 115274 531978
rect 115342 531922 115398 531978
rect 129250 597156 129306 597212
rect 129374 597156 129430 597212
rect 129498 597156 129554 597212
rect 129622 597156 129678 597212
rect 129250 597032 129306 597088
rect 129374 597032 129430 597088
rect 129498 597032 129554 597088
rect 129622 597032 129678 597088
rect 129250 596908 129306 596964
rect 129374 596908 129430 596964
rect 129498 596908 129554 596964
rect 129622 596908 129678 596964
rect 129250 596784 129306 596840
rect 129374 596784 129430 596840
rect 129498 596784 129554 596840
rect 129622 596784 129678 596840
rect 129250 580294 129306 580350
rect 129374 580294 129430 580350
rect 129498 580294 129554 580350
rect 129622 580294 129678 580350
rect 129250 580170 129306 580226
rect 129374 580170 129430 580226
rect 129498 580170 129554 580226
rect 129622 580170 129678 580226
rect 129250 580046 129306 580102
rect 129374 580046 129430 580102
rect 129498 580046 129554 580102
rect 129622 580046 129678 580102
rect 129250 579922 129306 579978
rect 129374 579922 129430 579978
rect 129498 579922 129554 579978
rect 129622 579922 129678 579978
rect 129250 562294 129306 562350
rect 129374 562294 129430 562350
rect 129498 562294 129554 562350
rect 129622 562294 129678 562350
rect 129250 562170 129306 562226
rect 129374 562170 129430 562226
rect 129498 562170 129554 562226
rect 129622 562170 129678 562226
rect 129250 562046 129306 562102
rect 129374 562046 129430 562102
rect 129498 562046 129554 562102
rect 129622 562046 129678 562102
rect 129250 561922 129306 561978
rect 129374 561922 129430 561978
rect 129498 561922 129554 561978
rect 129622 561922 129678 561978
rect 129250 544294 129306 544350
rect 129374 544294 129430 544350
rect 129498 544294 129554 544350
rect 129622 544294 129678 544350
rect 129250 544170 129306 544226
rect 129374 544170 129430 544226
rect 129498 544170 129554 544226
rect 129622 544170 129678 544226
rect 129250 544046 129306 544102
rect 129374 544046 129430 544102
rect 129498 544046 129554 544102
rect 129622 544046 129678 544102
rect 129250 543922 129306 543978
rect 129374 543922 129430 543978
rect 129498 543922 129554 543978
rect 129622 543922 129678 543978
rect 132970 598116 133026 598172
rect 133094 598116 133150 598172
rect 133218 598116 133274 598172
rect 133342 598116 133398 598172
rect 132970 597992 133026 598048
rect 133094 597992 133150 598048
rect 133218 597992 133274 598048
rect 133342 597992 133398 598048
rect 132970 597868 133026 597924
rect 133094 597868 133150 597924
rect 133218 597868 133274 597924
rect 133342 597868 133398 597924
rect 132970 597744 133026 597800
rect 133094 597744 133150 597800
rect 133218 597744 133274 597800
rect 133342 597744 133398 597800
rect 132970 586294 133026 586350
rect 133094 586294 133150 586350
rect 133218 586294 133274 586350
rect 133342 586294 133398 586350
rect 132970 586170 133026 586226
rect 133094 586170 133150 586226
rect 133218 586170 133274 586226
rect 133342 586170 133398 586226
rect 132970 586046 133026 586102
rect 133094 586046 133150 586102
rect 133218 586046 133274 586102
rect 133342 586046 133398 586102
rect 132970 585922 133026 585978
rect 133094 585922 133150 585978
rect 133218 585922 133274 585978
rect 133342 585922 133398 585978
rect 132970 568294 133026 568350
rect 133094 568294 133150 568350
rect 133218 568294 133274 568350
rect 133342 568294 133398 568350
rect 132970 568170 133026 568226
rect 133094 568170 133150 568226
rect 133218 568170 133274 568226
rect 133342 568170 133398 568226
rect 132970 568046 133026 568102
rect 133094 568046 133150 568102
rect 133218 568046 133274 568102
rect 133342 568046 133398 568102
rect 132970 567922 133026 567978
rect 133094 567922 133150 567978
rect 133218 567922 133274 567978
rect 133342 567922 133398 567978
rect 132970 550294 133026 550350
rect 133094 550294 133150 550350
rect 133218 550294 133274 550350
rect 133342 550294 133398 550350
rect 132970 550170 133026 550226
rect 133094 550170 133150 550226
rect 133218 550170 133274 550226
rect 133342 550170 133398 550226
rect 132970 550046 133026 550102
rect 133094 550046 133150 550102
rect 133218 550046 133274 550102
rect 133342 550046 133398 550102
rect 132970 549922 133026 549978
rect 133094 549922 133150 549978
rect 133218 549922 133274 549978
rect 133342 549922 133398 549978
rect 132970 532294 133026 532350
rect 133094 532294 133150 532350
rect 133218 532294 133274 532350
rect 133342 532294 133398 532350
rect 132970 532170 133026 532226
rect 133094 532170 133150 532226
rect 133218 532170 133274 532226
rect 133342 532170 133398 532226
rect 132970 532046 133026 532102
rect 133094 532046 133150 532102
rect 133218 532046 133274 532102
rect 133342 532046 133398 532102
rect 132970 531922 133026 531978
rect 133094 531922 133150 531978
rect 133218 531922 133274 531978
rect 133342 531922 133398 531978
rect 147250 597156 147306 597212
rect 147374 597156 147430 597212
rect 147498 597156 147554 597212
rect 147622 597156 147678 597212
rect 147250 597032 147306 597088
rect 147374 597032 147430 597088
rect 147498 597032 147554 597088
rect 147622 597032 147678 597088
rect 147250 596908 147306 596964
rect 147374 596908 147430 596964
rect 147498 596908 147554 596964
rect 147622 596908 147678 596964
rect 147250 596784 147306 596840
rect 147374 596784 147430 596840
rect 147498 596784 147554 596840
rect 147622 596784 147678 596840
rect 147250 580294 147306 580350
rect 147374 580294 147430 580350
rect 147498 580294 147554 580350
rect 147622 580294 147678 580350
rect 147250 580170 147306 580226
rect 147374 580170 147430 580226
rect 147498 580170 147554 580226
rect 147622 580170 147678 580226
rect 147250 580046 147306 580102
rect 147374 580046 147430 580102
rect 147498 580046 147554 580102
rect 147622 580046 147678 580102
rect 147250 579922 147306 579978
rect 147374 579922 147430 579978
rect 147498 579922 147554 579978
rect 147622 579922 147678 579978
rect 147250 562294 147306 562350
rect 147374 562294 147430 562350
rect 147498 562294 147554 562350
rect 147622 562294 147678 562350
rect 147250 562170 147306 562226
rect 147374 562170 147430 562226
rect 147498 562170 147554 562226
rect 147622 562170 147678 562226
rect 147250 562046 147306 562102
rect 147374 562046 147430 562102
rect 147498 562046 147554 562102
rect 147622 562046 147678 562102
rect 147250 561922 147306 561978
rect 147374 561922 147430 561978
rect 147498 561922 147554 561978
rect 147622 561922 147678 561978
rect 147250 544294 147306 544350
rect 147374 544294 147430 544350
rect 147498 544294 147554 544350
rect 147622 544294 147678 544350
rect 147250 544170 147306 544226
rect 147374 544170 147430 544226
rect 147498 544170 147554 544226
rect 147622 544170 147678 544226
rect 147250 544046 147306 544102
rect 147374 544046 147430 544102
rect 147498 544046 147554 544102
rect 147622 544046 147678 544102
rect 147250 543922 147306 543978
rect 147374 543922 147430 543978
rect 147498 543922 147554 543978
rect 147622 543922 147678 543978
rect 150970 598116 151026 598172
rect 151094 598116 151150 598172
rect 151218 598116 151274 598172
rect 151342 598116 151398 598172
rect 150970 597992 151026 598048
rect 151094 597992 151150 598048
rect 151218 597992 151274 598048
rect 151342 597992 151398 598048
rect 150970 597868 151026 597924
rect 151094 597868 151150 597924
rect 151218 597868 151274 597924
rect 151342 597868 151398 597924
rect 150970 597744 151026 597800
rect 151094 597744 151150 597800
rect 151218 597744 151274 597800
rect 151342 597744 151398 597800
rect 150970 586294 151026 586350
rect 151094 586294 151150 586350
rect 151218 586294 151274 586350
rect 151342 586294 151398 586350
rect 150970 586170 151026 586226
rect 151094 586170 151150 586226
rect 151218 586170 151274 586226
rect 151342 586170 151398 586226
rect 150970 586046 151026 586102
rect 151094 586046 151150 586102
rect 151218 586046 151274 586102
rect 151342 586046 151398 586102
rect 150970 585922 151026 585978
rect 151094 585922 151150 585978
rect 151218 585922 151274 585978
rect 151342 585922 151398 585978
rect 150970 568294 151026 568350
rect 151094 568294 151150 568350
rect 151218 568294 151274 568350
rect 151342 568294 151398 568350
rect 150970 568170 151026 568226
rect 151094 568170 151150 568226
rect 151218 568170 151274 568226
rect 151342 568170 151398 568226
rect 150970 568046 151026 568102
rect 151094 568046 151150 568102
rect 151218 568046 151274 568102
rect 151342 568046 151398 568102
rect 150970 567922 151026 567978
rect 151094 567922 151150 567978
rect 151218 567922 151274 567978
rect 151342 567922 151398 567978
rect 150970 550294 151026 550350
rect 151094 550294 151150 550350
rect 151218 550294 151274 550350
rect 151342 550294 151398 550350
rect 150970 550170 151026 550226
rect 151094 550170 151150 550226
rect 151218 550170 151274 550226
rect 151342 550170 151398 550226
rect 150970 550046 151026 550102
rect 151094 550046 151150 550102
rect 151218 550046 151274 550102
rect 151342 550046 151398 550102
rect 150970 549922 151026 549978
rect 151094 549922 151150 549978
rect 151218 549922 151274 549978
rect 151342 549922 151398 549978
rect 150970 532294 151026 532350
rect 151094 532294 151150 532350
rect 151218 532294 151274 532350
rect 151342 532294 151398 532350
rect 150970 532170 151026 532226
rect 151094 532170 151150 532226
rect 151218 532170 151274 532226
rect 151342 532170 151398 532226
rect 150970 532046 151026 532102
rect 151094 532046 151150 532102
rect 151218 532046 151274 532102
rect 151342 532046 151398 532102
rect 150970 531922 151026 531978
rect 151094 531922 151150 531978
rect 151218 531922 151274 531978
rect 151342 531922 151398 531978
rect 165250 597156 165306 597212
rect 165374 597156 165430 597212
rect 165498 597156 165554 597212
rect 165622 597156 165678 597212
rect 165250 597032 165306 597088
rect 165374 597032 165430 597088
rect 165498 597032 165554 597088
rect 165622 597032 165678 597088
rect 165250 596908 165306 596964
rect 165374 596908 165430 596964
rect 165498 596908 165554 596964
rect 165622 596908 165678 596964
rect 165250 596784 165306 596840
rect 165374 596784 165430 596840
rect 165498 596784 165554 596840
rect 165622 596784 165678 596840
rect 165250 580294 165306 580350
rect 165374 580294 165430 580350
rect 165498 580294 165554 580350
rect 165622 580294 165678 580350
rect 165250 580170 165306 580226
rect 165374 580170 165430 580226
rect 165498 580170 165554 580226
rect 165622 580170 165678 580226
rect 165250 580046 165306 580102
rect 165374 580046 165430 580102
rect 165498 580046 165554 580102
rect 165622 580046 165678 580102
rect 165250 579922 165306 579978
rect 165374 579922 165430 579978
rect 165498 579922 165554 579978
rect 165622 579922 165678 579978
rect 165250 562294 165306 562350
rect 165374 562294 165430 562350
rect 165498 562294 165554 562350
rect 165622 562294 165678 562350
rect 165250 562170 165306 562226
rect 165374 562170 165430 562226
rect 165498 562170 165554 562226
rect 165622 562170 165678 562226
rect 165250 562046 165306 562102
rect 165374 562046 165430 562102
rect 165498 562046 165554 562102
rect 165622 562046 165678 562102
rect 165250 561922 165306 561978
rect 165374 561922 165430 561978
rect 165498 561922 165554 561978
rect 165622 561922 165678 561978
rect 165250 544294 165306 544350
rect 165374 544294 165430 544350
rect 165498 544294 165554 544350
rect 165622 544294 165678 544350
rect 165250 544170 165306 544226
rect 165374 544170 165430 544226
rect 165498 544170 165554 544226
rect 165622 544170 165678 544226
rect 165250 544046 165306 544102
rect 165374 544046 165430 544102
rect 165498 544046 165554 544102
rect 165622 544046 165678 544102
rect 165250 543922 165306 543978
rect 165374 543922 165430 543978
rect 165498 543922 165554 543978
rect 165622 543922 165678 543978
rect 168970 598116 169026 598172
rect 169094 598116 169150 598172
rect 169218 598116 169274 598172
rect 169342 598116 169398 598172
rect 168970 597992 169026 598048
rect 169094 597992 169150 598048
rect 169218 597992 169274 598048
rect 169342 597992 169398 598048
rect 168970 597868 169026 597924
rect 169094 597868 169150 597924
rect 169218 597868 169274 597924
rect 169342 597868 169398 597924
rect 168970 597744 169026 597800
rect 169094 597744 169150 597800
rect 169218 597744 169274 597800
rect 169342 597744 169398 597800
rect 168970 586294 169026 586350
rect 169094 586294 169150 586350
rect 169218 586294 169274 586350
rect 169342 586294 169398 586350
rect 168970 586170 169026 586226
rect 169094 586170 169150 586226
rect 169218 586170 169274 586226
rect 169342 586170 169398 586226
rect 168970 586046 169026 586102
rect 169094 586046 169150 586102
rect 169218 586046 169274 586102
rect 169342 586046 169398 586102
rect 168970 585922 169026 585978
rect 169094 585922 169150 585978
rect 169218 585922 169274 585978
rect 169342 585922 169398 585978
rect 168970 568294 169026 568350
rect 169094 568294 169150 568350
rect 169218 568294 169274 568350
rect 169342 568294 169398 568350
rect 168970 568170 169026 568226
rect 169094 568170 169150 568226
rect 169218 568170 169274 568226
rect 169342 568170 169398 568226
rect 168970 568046 169026 568102
rect 169094 568046 169150 568102
rect 169218 568046 169274 568102
rect 169342 568046 169398 568102
rect 168970 567922 169026 567978
rect 169094 567922 169150 567978
rect 169218 567922 169274 567978
rect 169342 567922 169398 567978
rect 168970 550294 169026 550350
rect 169094 550294 169150 550350
rect 169218 550294 169274 550350
rect 169342 550294 169398 550350
rect 168970 550170 169026 550226
rect 169094 550170 169150 550226
rect 169218 550170 169274 550226
rect 169342 550170 169398 550226
rect 168970 550046 169026 550102
rect 169094 550046 169150 550102
rect 169218 550046 169274 550102
rect 169342 550046 169398 550102
rect 168970 549922 169026 549978
rect 169094 549922 169150 549978
rect 169218 549922 169274 549978
rect 169342 549922 169398 549978
rect 168970 532294 169026 532350
rect 169094 532294 169150 532350
rect 169218 532294 169274 532350
rect 169342 532294 169398 532350
rect 168970 532170 169026 532226
rect 169094 532170 169150 532226
rect 169218 532170 169274 532226
rect 169342 532170 169398 532226
rect 168970 532046 169026 532102
rect 169094 532046 169150 532102
rect 169218 532046 169274 532102
rect 169342 532046 169398 532102
rect 168970 531922 169026 531978
rect 169094 531922 169150 531978
rect 169218 531922 169274 531978
rect 169342 531922 169398 531978
rect 183250 597156 183306 597212
rect 183374 597156 183430 597212
rect 183498 597156 183554 597212
rect 183622 597156 183678 597212
rect 183250 597032 183306 597088
rect 183374 597032 183430 597088
rect 183498 597032 183554 597088
rect 183622 597032 183678 597088
rect 183250 596908 183306 596964
rect 183374 596908 183430 596964
rect 183498 596908 183554 596964
rect 183622 596908 183678 596964
rect 183250 596784 183306 596840
rect 183374 596784 183430 596840
rect 183498 596784 183554 596840
rect 183622 596784 183678 596840
rect 183250 580294 183306 580350
rect 183374 580294 183430 580350
rect 183498 580294 183554 580350
rect 183622 580294 183678 580350
rect 183250 580170 183306 580226
rect 183374 580170 183430 580226
rect 183498 580170 183554 580226
rect 183622 580170 183678 580226
rect 183250 580046 183306 580102
rect 183374 580046 183430 580102
rect 183498 580046 183554 580102
rect 183622 580046 183678 580102
rect 183250 579922 183306 579978
rect 183374 579922 183430 579978
rect 183498 579922 183554 579978
rect 183622 579922 183678 579978
rect 183250 562294 183306 562350
rect 183374 562294 183430 562350
rect 183498 562294 183554 562350
rect 183622 562294 183678 562350
rect 183250 562170 183306 562226
rect 183374 562170 183430 562226
rect 183498 562170 183554 562226
rect 183622 562170 183678 562226
rect 183250 562046 183306 562102
rect 183374 562046 183430 562102
rect 183498 562046 183554 562102
rect 183622 562046 183678 562102
rect 183250 561922 183306 561978
rect 183374 561922 183430 561978
rect 183498 561922 183554 561978
rect 183622 561922 183678 561978
rect 183250 544294 183306 544350
rect 183374 544294 183430 544350
rect 183498 544294 183554 544350
rect 183622 544294 183678 544350
rect 183250 544170 183306 544226
rect 183374 544170 183430 544226
rect 183498 544170 183554 544226
rect 183622 544170 183678 544226
rect 183250 544046 183306 544102
rect 183374 544046 183430 544102
rect 183498 544046 183554 544102
rect 183622 544046 183678 544102
rect 183250 543922 183306 543978
rect 183374 543922 183430 543978
rect 183498 543922 183554 543978
rect 183622 543922 183678 543978
rect 186970 598116 187026 598172
rect 187094 598116 187150 598172
rect 187218 598116 187274 598172
rect 187342 598116 187398 598172
rect 186970 597992 187026 598048
rect 187094 597992 187150 598048
rect 187218 597992 187274 598048
rect 187342 597992 187398 598048
rect 186970 597868 187026 597924
rect 187094 597868 187150 597924
rect 187218 597868 187274 597924
rect 187342 597868 187398 597924
rect 186970 597744 187026 597800
rect 187094 597744 187150 597800
rect 187218 597744 187274 597800
rect 187342 597744 187398 597800
rect 186970 586294 187026 586350
rect 187094 586294 187150 586350
rect 187218 586294 187274 586350
rect 187342 586294 187398 586350
rect 186970 586170 187026 586226
rect 187094 586170 187150 586226
rect 187218 586170 187274 586226
rect 187342 586170 187398 586226
rect 186970 586046 187026 586102
rect 187094 586046 187150 586102
rect 187218 586046 187274 586102
rect 187342 586046 187398 586102
rect 186970 585922 187026 585978
rect 187094 585922 187150 585978
rect 187218 585922 187274 585978
rect 187342 585922 187398 585978
rect 186970 568294 187026 568350
rect 187094 568294 187150 568350
rect 187218 568294 187274 568350
rect 187342 568294 187398 568350
rect 186970 568170 187026 568226
rect 187094 568170 187150 568226
rect 187218 568170 187274 568226
rect 187342 568170 187398 568226
rect 186970 568046 187026 568102
rect 187094 568046 187150 568102
rect 187218 568046 187274 568102
rect 187342 568046 187398 568102
rect 186970 567922 187026 567978
rect 187094 567922 187150 567978
rect 187218 567922 187274 567978
rect 187342 567922 187398 567978
rect 186970 550294 187026 550350
rect 187094 550294 187150 550350
rect 187218 550294 187274 550350
rect 187342 550294 187398 550350
rect 186970 550170 187026 550226
rect 187094 550170 187150 550226
rect 187218 550170 187274 550226
rect 187342 550170 187398 550226
rect 186970 550046 187026 550102
rect 187094 550046 187150 550102
rect 187218 550046 187274 550102
rect 187342 550046 187398 550102
rect 186970 549922 187026 549978
rect 187094 549922 187150 549978
rect 187218 549922 187274 549978
rect 187342 549922 187398 549978
rect 186970 532294 187026 532350
rect 187094 532294 187150 532350
rect 187218 532294 187274 532350
rect 187342 532294 187398 532350
rect 186970 532170 187026 532226
rect 187094 532170 187150 532226
rect 187218 532170 187274 532226
rect 187342 532170 187398 532226
rect 186970 532046 187026 532102
rect 187094 532046 187150 532102
rect 187218 532046 187274 532102
rect 187342 532046 187398 532102
rect 186970 531922 187026 531978
rect 187094 531922 187150 531978
rect 187218 531922 187274 531978
rect 187342 531922 187398 531978
rect 201250 597156 201306 597212
rect 201374 597156 201430 597212
rect 201498 597156 201554 597212
rect 201622 597156 201678 597212
rect 201250 597032 201306 597088
rect 201374 597032 201430 597088
rect 201498 597032 201554 597088
rect 201622 597032 201678 597088
rect 201250 596908 201306 596964
rect 201374 596908 201430 596964
rect 201498 596908 201554 596964
rect 201622 596908 201678 596964
rect 201250 596784 201306 596840
rect 201374 596784 201430 596840
rect 201498 596784 201554 596840
rect 201622 596784 201678 596840
rect 201250 580294 201306 580350
rect 201374 580294 201430 580350
rect 201498 580294 201554 580350
rect 201622 580294 201678 580350
rect 201250 580170 201306 580226
rect 201374 580170 201430 580226
rect 201498 580170 201554 580226
rect 201622 580170 201678 580226
rect 201250 580046 201306 580102
rect 201374 580046 201430 580102
rect 201498 580046 201554 580102
rect 201622 580046 201678 580102
rect 201250 579922 201306 579978
rect 201374 579922 201430 579978
rect 201498 579922 201554 579978
rect 201622 579922 201678 579978
rect 201250 562294 201306 562350
rect 201374 562294 201430 562350
rect 201498 562294 201554 562350
rect 201622 562294 201678 562350
rect 201250 562170 201306 562226
rect 201374 562170 201430 562226
rect 201498 562170 201554 562226
rect 201622 562170 201678 562226
rect 201250 562046 201306 562102
rect 201374 562046 201430 562102
rect 201498 562046 201554 562102
rect 201622 562046 201678 562102
rect 201250 561922 201306 561978
rect 201374 561922 201430 561978
rect 201498 561922 201554 561978
rect 201622 561922 201678 561978
rect 201250 544294 201306 544350
rect 201374 544294 201430 544350
rect 201498 544294 201554 544350
rect 201622 544294 201678 544350
rect 201250 544170 201306 544226
rect 201374 544170 201430 544226
rect 201498 544170 201554 544226
rect 201622 544170 201678 544226
rect 201250 544046 201306 544102
rect 201374 544046 201430 544102
rect 201498 544046 201554 544102
rect 201622 544046 201678 544102
rect 201250 543922 201306 543978
rect 201374 543922 201430 543978
rect 201498 543922 201554 543978
rect 201622 543922 201678 543978
rect 204970 598116 205026 598172
rect 205094 598116 205150 598172
rect 205218 598116 205274 598172
rect 205342 598116 205398 598172
rect 204970 597992 205026 598048
rect 205094 597992 205150 598048
rect 205218 597992 205274 598048
rect 205342 597992 205398 598048
rect 204970 597868 205026 597924
rect 205094 597868 205150 597924
rect 205218 597868 205274 597924
rect 205342 597868 205398 597924
rect 204970 597744 205026 597800
rect 205094 597744 205150 597800
rect 205218 597744 205274 597800
rect 205342 597744 205398 597800
rect 204970 586294 205026 586350
rect 205094 586294 205150 586350
rect 205218 586294 205274 586350
rect 205342 586294 205398 586350
rect 204970 586170 205026 586226
rect 205094 586170 205150 586226
rect 205218 586170 205274 586226
rect 205342 586170 205398 586226
rect 204970 586046 205026 586102
rect 205094 586046 205150 586102
rect 205218 586046 205274 586102
rect 205342 586046 205398 586102
rect 204970 585922 205026 585978
rect 205094 585922 205150 585978
rect 205218 585922 205274 585978
rect 205342 585922 205398 585978
rect 204970 568294 205026 568350
rect 205094 568294 205150 568350
rect 205218 568294 205274 568350
rect 205342 568294 205398 568350
rect 204970 568170 205026 568226
rect 205094 568170 205150 568226
rect 205218 568170 205274 568226
rect 205342 568170 205398 568226
rect 204970 568046 205026 568102
rect 205094 568046 205150 568102
rect 205218 568046 205274 568102
rect 205342 568046 205398 568102
rect 204970 567922 205026 567978
rect 205094 567922 205150 567978
rect 205218 567922 205274 567978
rect 205342 567922 205398 567978
rect 204970 550294 205026 550350
rect 205094 550294 205150 550350
rect 205218 550294 205274 550350
rect 205342 550294 205398 550350
rect 204970 550170 205026 550226
rect 205094 550170 205150 550226
rect 205218 550170 205274 550226
rect 205342 550170 205398 550226
rect 204970 550046 205026 550102
rect 205094 550046 205150 550102
rect 205218 550046 205274 550102
rect 205342 550046 205398 550102
rect 204970 549922 205026 549978
rect 205094 549922 205150 549978
rect 205218 549922 205274 549978
rect 205342 549922 205398 549978
rect 204970 532294 205026 532350
rect 205094 532294 205150 532350
rect 205218 532294 205274 532350
rect 205342 532294 205398 532350
rect 204970 532170 205026 532226
rect 205094 532170 205150 532226
rect 205218 532170 205274 532226
rect 205342 532170 205398 532226
rect 204970 532046 205026 532102
rect 205094 532046 205150 532102
rect 205218 532046 205274 532102
rect 205342 532046 205398 532102
rect 204970 531922 205026 531978
rect 205094 531922 205150 531978
rect 205218 531922 205274 531978
rect 205342 531922 205398 531978
rect 219250 597156 219306 597212
rect 219374 597156 219430 597212
rect 219498 597156 219554 597212
rect 219622 597156 219678 597212
rect 219250 597032 219306 597088
rect 219374 597032 219430 597088
rect 219498 597032 219554 597088
rect 219622 597032 219678 597088
rect 219250 596908 219306 596964
rect 219374 596908 219430 596964
rect 219498 596908 219554 596964
rect 219622 596908 219678 596964
rect 219250 596784 219306 596840
rect 219374 596784 219430 596840
rect 219498 596784 219554 596840
rect 219622 596784 219678 596840
rect 219250 580294 219306 580350
rect 219374 580294 219430 580350
rect 219498 580294 219554 580350
rect 219622 580294 219678 580350
rect 219250 580170 219306 580226
rect 219374 580170 219430 580226
rect 219498 580170 219554 580226
rect 219622 580170 219678 580226
rect 219250 580046 219306 580102
rect 219374 580046 219430 580102
rect 219498 580046 219554 580102
rect 219622 580046 219678 580102
rect 219250 579922 219306 579978
rect 219374 579922 219430 579978
rect 219498 579922 219554 579978
rect 219622 579922 219678 579978
rect 219250 562294 219306 562350
rect 219374 562294 219430 562350
rect 219498 562294 219554 562350
rect 219622 562294 219678 562350
rect 219250 562170 219306 562226
rect 219374 562170 219430 562226
rect 219498 562170 219554 562226
rect 219622 562170 219678 562226
rect 219250 562046 219306 562102
rect 219374 562046 219430 562102
rect 219498 562046 219554 562102
rect 219622 562046 219678 562102
rect 219250 561922 219306 561978
rect 219374 561922 219430 561978
rect 219498 561922 219554 561978
rect 219622 561922 219678 561978
rect 219250 544294 219306 544350
rect 219374 544294 219430 544350
rect 219498 544294 219554 544350
rect 219622 544294 219678 544350
rect 219250 544170 219306 544226
rect 219374 544170 219430 544226
rect 219498 544170 219554 544226
rect 219622 544170 219678 544226
rect 219250 544046 219306 544102
rect 219374 544046 219430 544102
rect 219498 544046 219554 544102
rect 219622 544046 219678 544102
rect 219250 543922 219306 543978
rect 219374 543922 219430 543978
rect 219498 543922 219554 543978
rect 219622 543922 219678 543978
rect 222970 598116 223026 598172
rect 223094 598116 223150 598172
rect 223218 598116 223274 598172
rect 223342 598116 223398 598172
rect 222970 597992 223026 598048
rect 223094 597992 223150 598048
rect 223218 597992 223274 598048
rect 223342 597992 223398 598048
rect 222970 597868 223026 597924
rect 223094 597868 223150 597924
rect 223218 597868 223274 597924
rect 223342 597868 223398 597924
rect 222970 597744 223026 597800
rect 223094 597744 223150 597800
rect 223218 597744 223274 597800
rect 223342 597744 223398 597800
rect 222970 586294 223026 586350
rect 223094 586294 223150 586350
rect 223218 586294 223274 586350
rect 223342 586294 223398 586350
rect 222970 586170 223026 586226
rect 223094 586170 223150 586226
rect 223218 586170 223274 586226
rect 223342 586170 223398 586226
rect 222970 586046 223026 586102
rect 223094 586046 223150 586102
rect 223218 586046 223274 586102
rect 223342 586046 223398 586102
rect 222970 585922 223026 585978
rect 223094 585922 223150 585978
rect 223218 585922 223274 585978
rect 223342 585922 223398 585978
rect 222970 568294 223026 568350
rect 223094 568294 223150 568350
rect 223218 568294 223274 568350
rect 223342 568294 223398 568350
rect 222970 568170 223026 568226
rect 223094 568170 223150 568226
rect 223218 568170 223274 568226
rect 223342 568170 223398 568226
rect 222970 568046 223026 568102
rect 223094 568046 223150 568102
rect 223218 568046 223274 568102
rect 223342 568046 223398 568102
rect 222970 567922 223026 567978
rect 223094 567922 223150 567978
rect 223218 567922 223274 567978
rect 223342 567922 223398 567978
rect 222970 550294 223026 550350
rect 223094 550294 223150 550350
rect 223218 550294 223274 550350
rect 223342 550294 223398 550350
rect 222970 550170 223026 550226
rect 223094 550170 223150 550226
rect 223218 550170 223274 550226
rect 223342 550170 223398 550226
rect 222970 550046 223026 550102
rect 223094 550046 223150 550102
rect 223218 550046 223274 550102
rect 223342 550046 223398 550102
rect 222970 549922 223026 549978
rect 223094 549922 223150 549978
rect 223218 549922 223274 549978
rect 223342 549922 223398 549978
rect 222970 532294 223026 532350
rect 223094 532294 223150 532350
rect 223218 532294 223274 532350
rect 223342 532294 223398 532350
rect 222970 532170 223026 532226
rect 223094 532170 223150 532226
rect 223218 532170 223274 532226
rect 223342 532170 223398 532226
rect 222970 532046 223026 532102
rect 223094 532046 223150 532102
rect 223218 532046 223274 532102
rect 223342 532046 223398 532102
rect 222970 531922 223026 531978
rect 223094 531922 223150 531978
rect 223218 531922 223274 531978
rect 223342 531922 223398 531978
rect 237250 597156 237306 597212
rect 237374 597156 237430 597212
rect 237498 597156 237554 597212
rect 237622 597156 237678 597212
rect 237250 597032 237306 597088
rect 237374 597032 237430 597088
rect 237498 597032 237554 597088
rect 237622 597032 237678 597088
rect 237250 596908 237306 596964
rect 237374 596908 237430 596964
rect 237498 596908 237554 596964
rect 237622 596908 237678 596964
rect 237250 596784 237306 596840
rect 237374 596784 237430 596840
rect 237498 596784 237554 596840
rect 237622 596784 237678 596840
rect 237250 580294 237306 580350
rect 237374 580294 237430 580350
rect 237498 580294 237554 580350
rect 237622 580294 237678 580350
rect 237250 580170 237306 580226
rect 237374 580170 237430 580226
rect 237498 580170 237554 580226
rect 237622 580170 237678 580226
rect 237250 580046 237306 580102
rect 237374 580046 237430 580102
rect 237498 580046 237554 580102
rect 237622 580046 237678 580102
rect 237250 579922 237306 579978
rect 237374 579922 237430 579978
rect 237498 579922 237554 579978
rect 237622 579922 237678 579978
rect 237250 562294 237306 562350
rect 237374 562294 237430 562350
rect 237498 562294 237554 562350
rect 237622 562294 237678 562350
rect 237250 562170 237306 562226
rect 237374 562170 237430 562226
rect 237498 562170 237554 562226
rect 237622 562170 237678 562226
rect 237250 562046 237306 562102
rect 237374 562046 237430 562102
rect 237498 562046 237554 562102
rect 237622 562046 237678 562102
rect 237250 561922 237306 561978
rect 237374 561922 237430 561978
rect 237498 561922 237554 561978
rect 237622 561922 237678 561978
rect 237250 544294 237306 544350
rect 237374 544294 237430 544350
rect 237498 544294 237554 544350
rect 237622 544294 237678 544350
rect 237250 544170 237306 544226
rect 237374 544170 237430 544226
rect 237498 544170 237554 544226
rect 237622 544170 237678 544226
rect 237250 544046 237306 544102
rect 237374 544046 237430 544102
rect 237498 544046 237554 544102
rect 237622 544046 237678 544102
rect 237250 543922 237306 543978
rect 237374 543922 237430 543978
rect 237498 543922 237554 543978
rect 237622 543922 237678 543978
rect 240970 598116 241026 598172
rect 241094 598116 241150 598172
rect 241218 598116 241274 598172
rect 241342 598116 241398 598172
rect 240970 597992 241026 598048
rect 241094 597992 241150 598048
rect 241218 597992 241274 598048
rect 241342 597992 241398 598048
rect 240970 597868 241026 597924
rect 241094 597868 241150 597924
rect 241218 597868 241274 597924
rect 241342 597868 241398 597924
rect 240970 597744 241026 597800
rect 241094 597744 241150 597800
rect 241218 597744 241274 597800
rect 241342 597744 241398 597800
rect 240970 586294 241026 586350
rect 241094 586294 241150 586350
rect 241218 586294 241274 586350
rect 241342 586294 241398 586350
rect 240970 586170 241026 586226
rect 241094 586170 241150 586226
rect 241218 586170 241274 586226
rect 241342 586170 241398 586226
rect 240970 586046 241026 586102
rect 241094 586046 241150 586102
rect 241218 586046 241274 586102
rect 241342 586046 241398 586102
rect 240970 585922 241026 585978
rect 241094 585922 241150 585978
rect 241218 585922 241274 585978
rect 241342 585922 241398 585978
rect 240970 568294 241026 568350
rect 241094 568294 241150 568350
rect 241218 568294 241274 568350
rect 241342 568294 241398 568350
rect 240970 568170 241026 568226
rect 241094 568170 241150 568226
rect 241218 568170 241274 568226
rect 241342 568170 241398 568226
rect 240970 568046 241026 568102
rect 241094 568046 241150 568102
rect 241218 568046 241274 568102
rect 241342 568046 241398 568102
rect 240970 567922 241026 567978
rect 241094 567922 241150 567978
rect 241218 567922 241274 567978
rect 241342 567922 241398 567978
rect 240970 550294 241026 550350
rect 241094 550294 241150 550350
rect 241218 550294 241274 550350
rect 241342 550294 241398 550350
rect 240970 550170 241026 550226
rect 241094 550170 241150 550226
rect 241218 550170 241274 550226
rect 241342 550170 241398 550226
rect 240970 550046 241026 550102
rect 241094 550046 241150 550102
rect 241218 550046 241274 550102
rect 241342 550046 241398 550102
rect 240970 549922 241026 549978
rect 241094 549922 241150 549978
rect 241218 549922 241274 549978
rect 241342 549922 241398 549978
rect 240970 532294 241026 532350
rect 241094 532294 241150 532350
rect 241218 532294 241274 532350
rect 241342 532294 241398 532350
rect 240970 532170 241026 532226
rect 241094 532170 241150 532226
rect 241218 532170 241274 532226
rect 241342 532170 241398 532226
rect 240970 532046 241026 532102
rect 241094 532046 241150 532102
rect 241218 532046 241274 532102
rect 241342 532046 241398 532102
rect 240970 531922 241026 531978
rect 241094 531922 241150 531978
rect 241218 531922 241274 531978
rect 241342 531922 241398 531978
rect 255250 597156 255306 597212
rect 255374 597156 255430 597212
rect 255498 597156 255554 597212
rect 255622 597156 255678 597212
rect 255250 597032 255306 597088
rect 255374 597032 255430 597088
rect 255498 597032 255554 597088
rect 255622 597032 255678 597088
rect 255250 596908 255306 596964
rect 255374 596908 255430 596964
rect 255498 596908 255554 596964
rect 255622 596908 255678 596964
rect 255250 596784 255306 596840
rect 255374 596784 255430 596840
rect 255498 596784 255554 596840
rect 255622 596784 255678 596840
rect 255250 580294 255306 580350
rect 255374 580294 255430 580350
rect 255498 580294 255554 580350
rect 255622 580294 255678 580350
rect 255250 580170 255306 580226
rect 255374 580170 255430 580226
rect 255498 580170 255554 580226
rect 255622 580170 255678 580226
rect 255250 580046 255306 580102
rect 255374 580046 255430 580102
rect 255498 580046 255554 580102
rect 255622 580046 255678 580102
rect 255250 579922 255306 579978
rect 255374 579922 255430 579978
rect 255498 579922 255554 579978
rect 255622 579922 255678 579978
rect 255250 562294 255306 562350
rect 255374 562294 255430 562350
rect 255498 562294 255554 562350
rect 255622 562294 255678 562350
rect 255250 562170 255306 562226
rect 255374 562170 255430 562226
rect 255498 562170 255554 562226
rect 255622 562170 255678 562226
rect 255250 562046 255306 562102
rect 255374 562046 255430 562102
rect 255498 562046 255554 562102
rect 255622 562046 255678 562102
rect 255250 561922 255306 561978
rect 255374 561922 255430 561978
rect 255498 561922 255554 561978
rect 255622 561922 255678 561978
rect 255250 544294 255306 544350
rect 255374 544294 255430 544350
rect 255498 544294 255554 544350
rect 255622 544294 255678 544350
rect 255250 544170 255306 544226
rect 255374 544170 255430 544226
rect 255498 544170 255554 544226
rect 255622 544170 255678 544226
rect 255250 544046 255306 544102
rect 255374 544046 255430 544102
rect 255498 544046 255554 544102
rect 255622 544046 255678 544102
rect 255250 543922 255306 543978
rect 255374 543922 255430 543978
rect 255498 543922 255554 543978
rect 255622 543922 255678 543978
rect 258970 598116 259026 598172
rect 259094 598116 259150 598172
rect 259218 598116 259274 598172
rect 259342 598116 259398 598172
rect 258970 597992 259026 598048
rect 259094 597992 259150 598048
rect 259218 597992 259274 598048
rect 259342 597992 259398 598048
rect 258970 597868 259026 597924
rect 259094 597868 259150 597924
rect 259218 597868 259274 597924
rect 259342 597868 259398 597924
rect 258970 597744 259026 597800
rect 259094 597744 259150 597800
rect 259218 597744 259274 597800
rect 259342 597744 259398 597800
rect 258970 586294 259026 586350
rect 259094 586294 259150 586350
rect 259218 586294 259274 586350
rect 259342 586294 259398 586350
rect 258970 586170 259026 586226
rect 259094 586170 259150 586226
rect 259218 586170 259274 586226
rect 259342 586170 259398 586226
rect 258970 586046 259026 586102
rect 259094 586046 259150 586102
rect 259218 586046 259274 586102
rect 259342 586046 259398 586102
rect 258970 585922 259026 585978
rect 259094 585922 259150 585978
rect 259218 585922 259274 585978
rect 259342 585922 259398 585978
rect 258970 568294 259026 568350
rect 259094 568294 259150 568350
rect 259218 568294 259274 568350
rect 259342 568294 259398 568350
rect 258970 568170 259026 568226
rect 259094 568170 259150 568226
rect 259218 568170 259274 568226
rect 259342 568170 259398 568226
rect 258970 568046 259026 568102
rect 259094 568046 259150 568102
rect 259218 568046 259274 568102
rect 259342 568046 259398 568102
rect 258970 567922 259026 567978
rect 259094 567922 259150 567978
rect 259218 567922 259274 567978
rect 259342 567922 259398 567978
rect 258970 550294 259026 550350
rect 259094 550294 259150 550350
rect 259218 550294 259274 550350
rect 259342 550294 259398 550350
rect 258970 550170 259026 550226
rect 259094 550170 259150 550226
rect 259218 550170 259274 550226
rect 259342 550170 259398 550226
rect 258970 550046 259026 550102
rect 259094 550046 259150 550102
rect 259218 550046 259274 550102
rect 259342 550046 259398 550102
rect 258970 549922 259026 549978
rect 259094 549922 259150 549978
rect 259218 549922 259274 549978
rect 259342 549922 259398 549978
rect 258970 532294 259026 532350
rect 259094 532294 259150 532350
rect 259218 532294 259274 532350
rect 259342 532294 259398 532350
rect 258970 532170 259026 532226
rect 259094 532170 259150 532226
rect 259218 532170 259274 532226
rect 259342 532170 259398 532226
rect 258970 532046 259026 532102
rect 259094 532046 259150 532102
rect 259218 532046 259274 532102
rect 259342 532046 259398 532102
rect 258970 531922 259026 531978
rect 259094 531922 259150 531978
rect 259218 531922 259274 531978
rect 259342 531922 259398 531978
rect 273250 597156 273306 597212
rect 273374 597156 273430 597212
rect 273498 597156 273554 597212
rect 273622 597156 273678 597212
rect 273250 597032 273306 597088
rect 273374 597032 273430 597088
rect 273498 597032 273554 597088
rect 273622 597032 273678 597088
rect 273250 596908 273306 596964
rect 273374 596908 273430 596964
rect 273498 596908 273554 596964
rect 273622 596908 273678 596964
rect 273250 596784 273306 596840
rect 273374 596784 273430 596840
rect 273498 596784 273554 596840
rect 273622 596784 273678 596840
rect 273250 580294 273306 580350
rect 273374 580294 273430 580350
rect 273498 580294 273554 580350
rect 273622 580294 273678 580350
rect 273250 580170 273306 580226
rect 273374 580170 273430 580226
rect 273498 580170 273554 580226
rect 273622 580170 273678 580226
rect 273250 580046 273306 580102
rect 273374 580046 273430 580102
rect 273498 580046 273554 580102
rect 273622 580046 273678 580102
rect 273250 579922 273306 579978
rect 273374 579922 273430 579978
rect 273498 579922 273554 579978
rect 273622 579922 273678 579978
rect 273250 562294 273306 562350
rect 273374 562294 273430 562350
rect 273498 562294 273554 562350
rect 273622 562294 273678 562350
rect 273250 562170 273306 562226
rect 273374 562170 273430 562226
rect 273498 562170 273554 562226
rect 273622 562170 273678 562226
rect 273250 562046 273306 562102
rect 273374 562046 273430 562102
rect 273498 562046 273554 562102
rect 273622 562046 273678 562102
rect 273250 561922 273306 561978
rect 273374 561922 273430 561978
rect 273498 561922 273554 561978
rect 273622 561922 273678 561978
rect 273250 544294 273306 544350
rect 273374 544294 273430 544350
rect 273498 544294 273554 544350
rect 273622 544294 273678 544350
rect 273250 544170 273306 544226
rect 273374 544170 273430 544226
rect 273498 544170 273554 544226
rect 273622 544170 273678 544226
rect 273250 544046 273306 544102
rect 273374 544046 273430 544102
rect 273498 544046 273554 544102
rect 273622 544046 273678 544102
rect 273250 543922 273306 543978
rect 273374 543922 273430 543978
rect 273498 543922 273554 543978
rect 273622 543922 273678 543978
rect 276970 598116 277026 598172
rect 277094 598116 277150 598172
rect 277218 598116 277274 598172
rect 277342 598116 277398 598172
rect 276970 597992 277026 598048
rect 277094 597992 277150 598048
rect 277218 597992 277274 598048
rect 277342 597992 277398 598048
rect 276970 597868 277026 597924
rect 277094 597868 277150 597924
rect 277218 597868 277274 597924
rect 277342 597868 277398 597924
rect 276970 597744 277026 597800
rect 277094 597744 277150 597800
rect 277218 597744 277274 597800
rect 277342 597744 277398 597800
rect 276970 586294 277026 586350
rect 277094 586294 277150 586350
rect 277218 586294 277274 586350
rect 277342 586294 277398 586350
rect 276970 586170 277026 586226
rect 277094 586170 277150 586226
rect 277218 586170 277274 586226
rect 277342 586170 277398 586226
rect 276970 586046 277026 586102
rect 277094 586046 277150 586102
rect 277218 586046 277274 586102
rect 277342 586046 277398 586102
rect 276970 585922 277026 585978
rect 277094 585922 277150 585978
rect 277218 585922 277274 585978
rect 277342 585922 277398 585978
rect 276970 568294 277026 568350
rect 277094 568294 277150 568350
rect 277218 568294 277274 568350
rect 277342 568294 277398 568350
rect 276970 568170 277026 568226
rect 277094 568170 277150 568226
rect 277218 568170 277274 568226
rect 277342 568170 277398 568226
rect 276970 568046 277026 568102
rect 277094 568046 277150 568102
rect 277218 568046 277274 568102
rect 277342 568046 277398 568102
rect 276970 567922 277026 567978
rect 277094 567922 277150 567978
rect 277218 567922 277274 567978
rect 277342 567922 277398 567978
rect 276970 550294 277026 550350
rect 277094 550294 277150 550350
rect 277218 550294 277274 550350
rect 277342 550294 277398 550350
rect 276970 550170 277026 550226
rect 277094 550170 277150 550226
rect 277218 550170 277274 550226
rect 277342 550170 277398 550226
rect 276970 550046 277026 550102
rect 277094 550046 277150 550102
rect 277218 550046 277274 550102
rect 277342 550046 277398 550102
rect 276970 549922 277026 549978
rect 277094 549922 277150 549978
rect 277218 549922 277274 549978
rect 277342 549922 277398 549978
rect 276970 532294 277026 532350
rect 277094 532294 277150 532350
rect 277218 532294 277274 532350
rect 277342 532294 277398 532350
rect 276970 532170 277026 532226
rect 277094 532170 277150 532226
rect 277218 532170 277274 532226
rect 277342 532170 277398 532226
rect 276970 532046 277026 532102
rect 277094 532046 277150 532102
rect 277218 532046 277274 532102
rect 277342 532046 277398 532102
rect 276970 531922 277026 531978
rect 277094 531922 277150 531978
rect 277218 531922 277274 531978
rect 277342 531922 277398 531978
rect 291250 597156 291306 597212
rect 291374 597156 291430 597212
rect 291498 597156 291554 597212
rect 291622 597156 291678 597212
rect 291250 597032 291306 597088
rect 291374 597032 291430 597088
rect 291498 597032 291554 597088
rect 291622 597032 291678 597088
rect 291250 596908 291306 596964
rect 291374 596908 291430 596964
rect 291498 596908 291554 596964
rect 291622 596908 291678 596964
rect 291250 596784 291306 596840
rect 291374 596784 291430 596840
rect 291498 596784 291554 596840
rect 291622 596784 291678 596840
rect 291250 580294 291306 580350
rect 291374 580294 291430 580350
rect 291498 580294 291554 580350
rect 291622 580294 291678 580350
rect 291250 580170 291306 580226
rect 291374 580170 291430 580226
rect 291498 580170 291554 580226
rect 291622 580170 291678 580226
rect 291250 580046 291306 580102
rect 291374 580046 291430 580102
rect 291498 580046 291554 580102
rect 291622 580046 291678 580102
rect 291250 579922 291306 579978
rect 291374 579922 291430 579978
rect 291498 579922 291554 579978
rect 291622 579922 291678 579978
rect 291250 562294 291306 562350
rect 291374 562294 291430 562350
rect 291498 562294 291554 562350
rect 291622 562294 291678 562350
rect 291250 562170 291306 562226
rect 291374 562170 291430 562226
rect 291498 562170 291554 562226
rect 291622 562170 291678 562226
rect 291250 562046 291306 562102
rect 291374 562046 291430 562102
rect 291498 562046 291554 562102
rect 291622 562046 291678 562102
rect 291250 561922 291306 561978
rect 291374 561922 291430 561978
rect 291498 561922 291554 561978
rect 291622 561922 291678 561978
rect 291250 544294 291306 544350
rect 291374 544294 291430 544350
rect 291498 544294 291554 544350
rect 291622 544294 291678 544350
rect 291250 544170 291306 544226
rect 291374 544170 291430 544226
rect 291498 544170 291554 544226
rect 291622 544170 291678 544226
rect 291250 544046 291306 544102
rect 291374 544046 291430 544102
rect 291498 544046 291554 544102
rect 291622 544046 291678 544102
rect 291250 543922 291306 543978
rect 291374 543922 291430 543978
rect 291498 543922 291554 543978
rect 291622 543922 291678 543978
rect 294970 598116 295026 598172
rect 295094 598116 295150 598172
rect 295218 598116 295274 598172
rect 295342 598116 295398 598172
rect 294970 597992 295026 598048
rect 295094 597992 295150 598048
rect 295218 597992 295274 598048
rect 295342 597992 295398 598048
rect 294970 597868 295026 597924
rect 295094 597868 295150 597924
rect 295218 597868 295274 597924
rect 295342 597868 295398 597924
rect 294970 597744 295026 597800
rect 295094 597744 295150 597800
rect 295218 597744 295274 597800
rect 295342 597744 295398 597800
rect 294970 586294 295026 586350
rect 295094 586294 295150 586350
rect 295218 586294 295274 586350
rect 295342 586294 295398 586350
rect 294970 586170 295026 586226
rect 295094 586170 295150 586226
rect 295218 586170 295274 586226
rect 295342 586170 295398 586226
rect 294970 586046 295026 586102
rect 295094 586046 295150 586102
rect 295218 586046 295274 586102
rect 295342 586046 295398 586102
rect 294970 585922 295026 585978
rect 295094 585922 295150 585978
rect 295218 585922 295274 585978
rect 295342 585922 295398 585978
rect 294970 568294 295026 568350
rect 295094 568294 295150 568350
rect 295218 568294 295274 568350
rect 295342 568294 295398 568350
rect 294970 568170 295026 568226
rect 295094 568170 295150 568226
rect 295218 568170 295274 568226
rect 295342 568170 295398 568226
rect 294970 568046 295026 568102
rect 295094 568046 295150 568102
rect 295218 568046 295274 568102
rect 295342 568046 295398 568102
rect 294970 567922 295026 567978
rect 295094 567922 295150 567978
rect 295218 567922 295274 567978
rect 295342 567922 295398 567978
rect 294970 550294 295026 550350
rect 295094 550294 295150 550350
rect 295218 550294 295274 550350
rect 295342 550294 295398 550350
rect 294970 550170 295026 550226
rect 295094 550170 295150 550226
rect 295218 550170 295274 550226
rect 295342 550170 295398 550226
rect 294970 550046 295026 550102
rect 295094 550046 295150 550102
rect 295218 550046 295274 550102
rect 295342 550046 295398 550102
rect 294970 549922 295026 549978
rect 295094 549922 295150 549978
rect 295218 549922 295274 549978
rect 295342 549922 295398 549978
rect 294970 532294 295026 532350
rect 295094 532294 295150 532350
rect 295218 532294 295274 532350
rect 295342 532294 295398 532350
rect 294970 532170 295026 532226
rect 295094 532170 295150 532226
rect 295218 532170 295274 532226
rect 295342 532170 295398 532226
rect 294970 532046 295026 532102
rect 295094 532046 295150 532102
rect 295218 532046 295274 532102
rect 295342 532046 295398 532102
rect 294970 531922 295026 531978
rect 295094 531922 295150 531978
rect 295218 531922 295274 531978
rect 295342 531922 295398 531978
rect 309250 597156 309306 597212
rect 309374 597156 309430 597212
rect 309498 597156 309554 597212
rect 309622 597156 309678 597212
rect 309250 597032 309306 597088
rect 309374 597032 309430 597088
rect 309498 597032 309554 597088
rect 309622 597032 309678 597088
rect 309250 596908 309306 596964
rect 309374 596908 309430 596964
rect 309498 596908 309554 596964
rect 309622 596908 309678 596964
rect 309250 596784 309306 596840
rect 309374 596784 309430 596840
rect 309498 596784 309554 596840
rect 309622 596784 309678 596840
rect 309250 580294 309306 580350
rect 309374 580294 309430 580350
rect 309498 580294 309554 580350
rect 309622 580294 309678 580350
rect 309250 580170 309306 580226
rect 309374 580170 309430 580226
rect 309498 580170 309554 580226
rect 309622 580170 309678 580226
rect 309250 580046 309306 580102
rect 309374 580046 309430 580102
rect 309498 580046 309554 580102
rect 309622 580046 309678 580102
rect 309250 579922 309306 579978
rect 309374 579922 309430 579978
rect 309498 579922 309554 579978
rect 309622 579922 309678 579978
rect 309250 562294 309306 562350
rect 309374 562294 309430 562350
rect 309498 562294 309554 562350
rect 309622 562294 309678 562350
rect 309250 562170 309306 562226
rect 309374 562170 309430 562226
rect 309498 562170 309554 562226
rect 309622 562170 309678 562226
rect 309250 562046 309306 562102
rect 309374 562046 309430 562102
rect 309498 562046 309554 562102
rect 309622 562046 309678 562102
rect 309250 561922 309306 561978
rect 309374 561922 309430 561978
rect 309498 561922 309554 561978
rect 309622 561922 309678 561978
rect 309250 544294 309306 544350
rect 309374 544294 309430 544350
rect 309498 544294 309554 544350
rect 309622 544294 309678 544350
rect 309250 544170 309306 544226
rect 309374 544170 309430 544226
rect 309498 544170 309554 544226
rect 309622 544170 309678 544226
rect 309250 544046 309306 544102
rect 309374 544046 309430 544102
rect 309498 544046 309554 544102
rect 309622 544046 309678 544102
rect 309250 543922 309306 543978
rect 309374 543922 309430 543978
rect 309498 543922 309554 543978
rect 309622 543922 309678 543978
rect 312970 598116 313026 598172
rect 313094 598116 313150 598172
rect 313218 598116 313274 598172
rect 313342 598116 313398 598172
rect 312970 597992 313026 598048
rect 313094 597992 313150 598048
rect 313218 597992 313274 598048
rect 313342 597992 313398 598048
rect 312970 597868 313026 597924
rect 313094 597868 313150 597924
rect 313218 597868 313274 597924
rect 313342 597868 313398 597924
rect 312970 597744 313026 597800
rect 313094 597744 313150 597800
rect 313218 597744 313274 597800
rect 313342 597744 313398 597800
rect 312970 586294 313026 586350
rect 313094 586294 313150 586350
rect 313218 586294 313274 586350
rect 313342 586294 313398 586350
rect 312970 586170 313026 586226
rect 313094 586170 313150 586226
rect 313218 586170 313274 586226
rect 313342 586170 313398 586226
rect 312970 586046 313026 586102
rect 313094 586046 313150 586102
rect 313218 586046 313274 586102
rect 313342 586046 313398 586102
rect 312970 585922 313026 585978
rect 313094 585922 313150 585978
rect 313218 585922 313274 585978
rect 313342 585922 313398 585978
rect 312970 568294 313026 568350
rect 313094 568294 313150 568350
rect 313218 568294 313274 568350
rect 313342 568294 313398 568350
rect 312970 568170 313026 568226
rect 313094 568170 313150 568226
rect 313218 568170 313274 568226
rect 313342 568170 313398 568226
rect 312970 568046 313026 568102
rect 313094 568046 313150 568102
rect 313218 568046 313274 568102
rect 313342 568046 313398 568102
rect 312970 567922 313026 567978
rect 313094 567922 313150 567978
rect 313218 567922 313274 567978
rect 313342 567922 313398 567978
rect 312970 550294 313026 550350
rect 313094 550294 313150 550350
rect 313218 550294 313274 550350
rect 313342 550294 313398 550350
rect 312970 550170 313026 550226
rect 313094 550170 313150 550226
rect 313218 550170 313274 550226
rect 313342 550170 313398 550226
rect 312970 550046 313026 550102
rect 313094 550046 313150 550102
rect 313218 550046 313274 550102
rect 313342 550046 313398 550102
rect 312970 549922 313026 549978
rect 313094 549922 313150 549978
rect 313218 549922 313274 549978
rect 313342 549922 313398 549978
rect 312970 532294 313026 532350
rect 313094 532294 313150 532350
rect 313218 532294 313274 532350
rect 313342 532294 313398 532350
rect 312970 532170 313026 532226
rect 313094 532170 313150 532226
rect 313218 532170 313274 532226
rect 313342 532170 313398 532226
rect 312970 532046 313026 532102
rect 313094 532046 313150 532102
rect 313218 532046 313274 532102
rect 313342 532046 313398 532102
rect 312970 531922 313026 531978
rect 313094 531922 313150 531978
rect 313218 531922 313274 531978
rect 313342 531922 313398 531978
rect 327250 597156 327306 597212
rect 327374 597156 327430 597212
rect 327498 597156 327554 597212
rect 327622 597156 327678 597212
rect 327250 597032 327306 597088
rect 327374 597032 327430 597088
rect 327498 597032 327554 597088
rect 327622 597032 327678 597088
rect 327250 596908 327306 596964
rect 327374 596908 327430 596964
rect 327498 596908 327554 596964
rect 327622 596908 327678 596964
rect 327250 596784 327306 596840
rect 327374 596784 327430 596840
rect 327498 596784 327554 596840
rect 327622 596784 327678 596840
rect 327250 580294 327306 580350
rect 327374 580294 327430 580350
rect 327498 580294 327554 580350
rect 327622 580294 327678 580350
rect 327250 580170 327306 580226
rect 327374 580170 327430 580226
rect 327498 580170 327554 580226
rect 327622 580170 327678 580226
rect 327250 580046 327306 580102
rect 327374 580046 327430 580102
rect 327498 580046 327554 580102
rect 327622 580046 327678 580102
rect 327250 579922 327306 579978
rect 327374 579922 327430 579978
rect 327498 579922 327554 579978
rect 327622 579922 327678 579978
rect 327250 562294 327306 562350
rect 327374 562294 327430 562350
rect 327498 562294 327554 562350
rect 327622 562294 327678 562350
rect 327250 562170 327306 562226
rect 327374 562170 327430 562226
rect 327498 562170 327554 562226
rect 327622 562170 327678 562226
rect 327250 562046 327306 562102
rect 327374 562046 327430 562102
rect 327498 562046 327554 562102
rect 327622 562046 327678 562102
rect 327250 561922 327306 561978
rect 327374 561922 327430 561978
rect 327498 561922 327554 561978
rect 327622 561922 327678 561978
rect 327250 544294 327306 544350
rect 327374 544294 327430 544350
rect 327498 544294 327554 544350
rect 327622 544294 327678 544350
rect 327250 544170 327306 544226
rect 327374 544170 327430 544226
rect 327498 544170 327554 544226
rect 327622 544170 327678 544226
rect 327250 544046 327306 544102
rect 327374 544046 327430 544102
rect 327498 544046 327554 544102
rect 327622 544046 327678 544102
rect 327250 543922 327306 543978
rect 327374 543922 327430 543978
rect 327498 543922 327554 543978
rect 327622 543922 327678 543978
rect 330970 598116 331026 598172
rect 331094 598116 331150 598172
rect 331218 598116 331274 598172
rect 331342 598116 331398 598172
rect 330970 597992 331026 598048
rect 331094 597992 331150 598048
rect 331218 597992 331274 598048
rect 331342 597992 331398 598048
rect 330970 597868 331026 597924
rect 331094 597868 331150 597924
rect 331218 597868 331274 597924
rect 331342 597868 331398 597924
rect 330970 597744 331026 597800
rect 331094 597744 331150 597800
rect 331218 597744 331274 597800
rect 331342 597744 331398 597800
rect 330970 586294 331026 586350
rect 331094 586294 331150 586350
rect 331218 586294 331274 586350
rect 331342 586294 331398 586350
rect 330970 586170 331026 586226
rect 331094 586170 331150 586226
rect 331218 586170 331274 586226
rect 331342 586170 331398 586226
rect 330970 586046 331026 586102
rect 331094 586046 331150 586102
rect 331218 586046 331274 586102
rect 331342 586046 331398 586102
rect 330970 585922 331026 585978
rect 331094 585922 331150 585978
rect 331218 585922 331274 585978
rect 331342 585922 331398 585978
rect 330970 568294 331026 568350
rect 331094 568294 331150 568350
rect 331218 568294 331274 568350
rect 331342 568294 331398 568350
rect 330970 568170 331026 568226
rect 331094 568170 331150 568226
rect 331218 568170 331274 568226
rect 331342 568170 331398 568226
rect 330970 568046 331026 568102
rect 331094 568046 331150 568102
rect 331218 568046 331274 568102
rect 331342 568046 331398 568102
rect 330970 567922 331026 567978
rect 331094 567922 331150 567978
rect 331218 567922 331274 567978
rect 331342 567922 331398 567978
rect 330970 550294 331026 550350
rect 331094 550294 331150 550350
rect 331218 550294 331274 550350
rect 331342 550294 331398 550350
rect 330970 550170 331026 550226
rect 331094 550170 331150 550226
rect 331218 550170 331274 550226
rect 331342 550170 331398 550226
rect 330970 550046 331026 550102
rect 331094 550046 331150 550102
rect 331218 550046 331274 550102
rect 331342 550046 331398 550102
rect 330970 549922 331026 549978
rect 331094 549922 331150 549978
rect 331218 549922 331274 549978
rect 331342 549922 331398 549978
rect 330970 532294 331026 532350
rect 331094 532294 331150 532350
rect 331218 532294 331274 532350
rect 331342 532294 331398 532350
rect 330970 532170 331026 532226
rect 331094 532170 331150 532226
rect 331218 532170 331274 532226
rect 331342 532170 331398 532226
rect 330970 532046 331026 532102
rect 331094 532046 331150 532102
rect 331218 532046 331274 532102
rect 331342 532046 331398 532102
rect 330970 531922 331026 531978
rect 331094 531922 331150 531978
rect 331218 531922 331274 531978
rect 331342 531922 331398 531978
rect 345250 597156 345306 597212
rect 345374 597156 345430 597212
rect 345498 597156 345554 597212
rect 345622 597156 345678 597212
rect 345250 597032 345306 597088
rect 345374 597032 345430 597088
rect 345498 597032 345554 597088
rect 345622 597032 345678 597088
rect 345250 596908 345306 596964
rect 345374 596908 345430 596964
rect 345498 596908 345554 596964
rect 345622 596908 345678 596964
rect 345250 596784 345306 596840
rect 345374 596784 345430 596840
rect 345498 596784 345554 596840
rect 345622 596784 345678 596840
rect 345250 580294 345306 580350
rect 345374 580294 345430 580350
rect 345498 580294 345554 580350
rect 345622 580294 345678 580350
rect 345250 580170 345306 580226
rect 345374 580170 345430 580226
rect 345498 580170 345554 580226
rect 345622 580170 345678 580226
rect 345250 580046 345306 580102
rect 345374 580046 345430 580102
rect 345498 580046 345554 580102
rect 345622 580046 345678 580102
rect 345250 579922 345306 579978
rect 345374 579922 345430 579978
rect 345498 579922 345554 579978
rect 345622 579922 345678 579978
rect 345250 562294 345306 562350
rect 345374 562294 345430 562350
rect 345498 562294 345554 562350
rect 345622 562294 345678 562350
rect 345250 562170 345306 562226
rect 345374 562170 345430 562226
rect 345498 562170 345554 562226
rect 345622 562170 345678 562226
rect 345250 562046 345306 562102
rect 345374 562046 345430 562102
rect 345498 562046 345554 562102
rect 345622 562046 345678 562102
rect 345250 561922 345306 561978
rect 345374 561922 345430 561978
rect 345498 561922 345554 561978
rect 345622 561922 345678 561978
rect 345250 544294 345306 544350
rect 345374 544294 345430 544350
rect 345498 544294 345554 544350
rect 345622 544294 345678 544350
rect 345250 544170 345306 544226
rect 345374 544170 345430 544226
rect 345498 544170 345554 544226
rect 345622 544170 345678 544226
rect 345250 544046 345306 544102
rect 345374 544046 345430 544102
rect 345498 544046 345554 544102
rect 345622 544046 345678 544102
rect 345250 543922 345306 543978
rect 345374 543922 345430 543978
rect 345498 543922 345554 543978
rect 345622 543922 345678 543978
rect 348970 598116 349026 598172
rect 349094 598116 349150 598172
rect 349218 598116 349274 598172
rect 349342 598116 349398 598172
rect 348970 597992 349026 598048
rect 349094 597992 349150 598048
rect 349218 597992 349274 598048
rect 349342 597992 349398 598048
rect 348970 597868 349026 597924
rect 349094 597868 349150 597924
rect 349218 597868 349274 597924
rect 349342 597868 349398 597924
rect 348970 597744 349026 597800
rect 349094 597744 349150 597800
rect 349218 597744 349274 597800
rect 349342 597744 349398 597800
rect 348970 586294 349026 586350
rect 349094 586294 349150 586350
rect 349218 586294 349274 586350
rect 349342 586294 349398 586350
rect 348970 586170 349026 586226
rect 349094 586170 349150 586226
rect 349218 586170 349274 586226
rect 349342 586170 349398 586226
rect 348970 586046 349026 586102
rect 349094 586046 349150 586102
rect 349218 586046 349274 586102
rect 349342 586046 349398 586102
rect 348970 585922 349026 585978
rect 349094 585922 349150 585978
rect 349218 585922 349274 585978
rect 349342 585922 349398 585978
rect 348970 568294 349026 568350
rect 349094 568294 349150 568350
rect 349218 568294 349274 568350
rect 349342 568294 349398 568350
rect 348970 568170 349026 568226
rect 349094 568170 349150 568226
rect 349218 568170 349274 568226
rect 349342 568170 349398 568226
rect 348970 568046 349026 568102
rect 349094 568046 349150 568102
rect 349218 568046 349274 568102
rect 349342 568046 349398 568102
rect 348970 567922 349026 567978
rect 349094 567922 349150 567978
rect 349218 567922 349274 567978
rect 349342 567922 349398 567978
rect 348970 550294 349026 550350
rect 349094 550294 349150 550350
rect 349218 550294 349274 550350
rect 349342 550294 349398 550350
rect 348970 550170 349026 550226
rect 349094 550170 349150 550226
rect 349218 550170 349274 550226
rect 349342 550170 349398 550226
rect 348970 550046 349026 550102
rect 349094 550046 349150 550102
rect 349218 550046 349274 550102
rect 349342 550046 349398 550102
rect 348970 549922 349026 549978
rect 349094 549922 349150 549978
rect 349218 549922 349274 549978
rect 349342 549922 349398 549978
rect 348970 532294 349026 532350
rect 349094 532294 349150 532350
rect 349218 532294 349274 532350
rect 349342 532294 349398 532350
rect 348970 532170 349026 532226
rect 349094 532170 349150 532226
rect 349218 532170 349274 532226
rect 349342 532170 349398 532226
rect 348970 532046 349026 532102
rect 349094 532046 349150 532102
rect 349218 532046 349274 532102
rect 349342 532046 349398 532102
rect 348970 531922 349026 531978
rect 349094 531922 349150 531978
rect 349218 531922 349274 531978
rect 349342 531922 349398 531978
rect 363250 597156 363306 597212
rect 363374 597156 363430 597212
rect 363498 597156 363554 597212
rect 363622 597156 363678 597212
rect 363250 597032 363306 597088
rect 363374 597032 363430 597088
rect 363498 597032 363554 597088
rect 363622 597032 363678 597088
rect 363250 596908 363306 596964
rect 363374 596908 363430 596964
rect 363498 596908 363554 596964
rect 363622 596908 363678 596964
rect 363250 596784 363306 596840
rect 363374 596784 363430 596840
rect 363498 596784 363554 596840
rect 363622 596784 363678 596840
rect 363250 580294 363306 580350
rect 363374 580294 363430 580350
rect 363498 580294 363554 580350
rect 363622 580294 363678 580350
rect 363250 580170 363306 580226
rect 363374 580170 363430 580226
rect 363498 580170 363554 580226
rect 363622 580170 363678 580226
rect 363250 580046 363306 580102
rect 363374 580046 363430 580102
rect 363498 580046 363554 580102
rect 363622 580046 363678 580102
rect 363250 579922 363306 579978
rect 363374 579922 363430 579978
rect 363498 579922 363554 579978
rect 363622 579922 363678 579978
rect 363250 562294 363306 562350
rect 363374 562294 363430 562350
rect 363498 562294 363554 562350
rect 363622 562294 363678 562350
rect 363250 562170 363306 562226
rect 363374 562170 363430 562226
rect 363498 562170 363554 562226
rect 363622 562170 363678 562226
rect 363250 562046 363306 562102
rect 363374 562046 363430 562102
rect 363498 562046 363554 562102
rect 363622 562046 363678 562102
rect 363250 561922 363306 561978
rect 363374 561922 363430 561978
rect 363498 561922 363554 561978
rect 363622 561922 363678 561978
rect 363250 544294 363306 544350
rect 363374 544294 363430 544350
rect 363498 544294 363554 544350
rect 363622 544294 363678 544350
rect 363250 544170 363306 544226
rect 363374 544170 363430 544226
rect 363498 544170 363554 544226
rect 363622 544170 363678 544226
rect 363250 544046 363306 544102
rect 363374 544046 363430 544102
rect 363498 544046 363554 544102
rect 363622 544046 363678 544102
rect 363250 543922 363306 543978
rect 363374 543922 363430 543978
rect 363498 543922 363554 543978
rect 363622 543922 363678 543978
rect 366970 598116 367026 598172
rect 367094 598116 367150 598172
rect 367218 598116 367274 598172
rect 367342 598116 367398 598172
rect 366970 597992 367026 598048
rect 367094 597992 367150 598048
rect 367218 597992 367274 598048
rect 367342 597992 367398 598048
rect 366970 597868 367026 597924
rect 367094 597868 367150 597924
rect 367218 597868 367274 597924
rect 367342 597868 367398 597924
rect 366970 597744 367026 597800
rect 367094 597744 367150 597800
rect 367218 597744 367274 597800
rect 367342 597744 367398 597800
rect 366970 586294 367026 586350
rect 367094 586294 367150 586350
rect 367218 586294 367274 586350
rect 367342 586294 367398 586350
rect 366970 586170 367026 586226
rect 367094 586170 367150 586226
rect 367218 586170 367274 586226
rect 367342 586170 367398 586226
rect 366970 586046 367026 586102
rect 367094 586046 367150 586102
rect 367218 586046 367274 586102
rect 367342 586046 367398 586102
rect 366970 585922 367026 585978
rect 367094 585922 367150 585978
rect 367218 585922 367274 585978
rect 367342 585922 367398 585978
rect 366970 568294 367026 568350
rect 367094 568294 367150 568350
rect 367218 568294 367274 568350
rect 367342 568294 367398 568350
rect 366970 568170 367026 568226
rect 367094 568170 367150 568226
rect 367218 568170 367274 568226
rect 367342 568170 367398 568226
rect 366970 568046 367026 568102
rect 367094 568046 367150 568102
rect 367218 568046 367274 568102
rect 367342 568046 367398 568102
rect 366970 567922 367026 567978
rect 367094 567922 367150 567978
rect 367218 567922 367274 567978
rect 367342 567922 367398 567978
rect 366970 550294 367026 550350
rect 367094 550294 367150 550350
rect 367218 550294 367274 550350
rect 367342 550294 367398 550350
rect 366970 550170 367026 550226
rect 367094 550170 367150 550226
rect 367218 550170 367274 550226
rect 367342 550170 367398 550226
rect 366970 550046 367026 550102
rect 367094 550046 367150 550102
rect 367218 550046 367274 550102
rect 367342 550046 367398 550102
rect 366970 549922 367026 549978
rect 367094 549922 367150 549978
rect 367218 549922 367274 549978
rect 367342 549922 367398 549978
rect 366970 532294 367026 532350
rect 367094 532294 367150 532350
rect 367218 532294 367274 532350
rect 367342 532294 367398 532350
rect 366970 532170 367026 532226
rect 367094 532170 367150 532226
rect 367218 532170 367274 532226
rect 367342 532170 367398 532226
rect 366970 532046 367026 532102
rect 367094 532046 367150 532102
rect 367218 532046 367274 532102
rect 367342 532046 367398 532102
rect 366970 531922 367026 531978
rect 367094 531922 367150 531978
rect 367218 531922 367274 531978
rect 367342 531922 367398 531978
rect 381250 597156 381306 597212
rect 381374 597156 381430 597212
rect 381498 597156 381554 597212
rect 381622 597156 381678 597212
rect 381250 597032 381306 597088
rect 381374 597032 381430 597088
rect 381498 597032 381554 597088
rect 381622 597032 381678 597088
rect 381250 596908 381306 596964
rect 381374 596908 381430 596964
rect 381498 596908 381554 596964
rect 381622 596908 381678 596964
rect 381250 596784 381306 596840
rect 381374 596784 381430 596840
rect 381498 596784 381554 596840
rect 381622 596784 381678 596840
rect 381250 580294 381306 580350
rect 381374 580294 381430 580350
rect 381498 580294 381554 580350
rect 381622 580294 381678 580350
rect 381250 580170 381306 580226
rect 381374 580170 381430 580226
rect 381498 580170 381554 580226
rect 381622 580170 381678 580226
rect 381250 580046 381306 580102
rect 381374 580046 381430 580102
rect 381498 580046 381554 580102
rect 381622 580046 381678 580102
rect 381250 579922 381306 579978
rect 381374 579922 381430 579978
rect 381498 579922 381554 579978
rect 381622 579922 381678 579978
rect 381250 562294 381306 562350
rect 381374 562294 381430 562350
rect 381498 562294 381554 562350
rect 381622 562294 381678 562350
rect 381250 562170 381306 562226
rect 381374 562170 381430 562226
rect 381498 562170 381554 562226
rect 381622 562170 381678 562226
rect 381250 562046 381306 562102
rect 381374 562046 381430 562102
rect 381498 562046 381554 562102
rect 381622 562046 381678 562102
rect 381250 561922 381306 561978
rect 381374 561922 381430 561978
rect 381498 561922 381554 561978
rect 381622 561922 381678 561978
rect 381250 544294 381306 544350
rect 381374 544294 381430 544350
rect 381498 544294 381554 544350
rect 381622 544294 381678 544350
rect 381250 544170 381306 544226
rect 381374 544170 381430 544226
rect 381498 544170 381554 544226
rect 381622 544170 381678 544226
rect 381250 544046 381306 544102
rect 381374 544046 381430 544102
rect 381498 544046 381554 544102
rect 381622 544046 381678 544102
rect 381250 543922 381306 543978
rect 381374 543922 381430 543978
rect 381498 543922 381554 543978
rect 381622 543922 381678 543978
rect 384970 598116 385026 598172
rect 385094 598116 385150 598172
rect 385218 598116 385274 598172
rect 385342 598116 385398 598172
rect 384970 597992 385026 598048
rect 385094 597992 385150 598048
rect 385218 597992 385274 598048
rect 385342 597992 385398 598048
rect 384970 597868 385026 597924
rect 385094 597868 385150 597924
rect 385218 597868 385274 597924
rect 385342 597868 385398 597924
rect 384970 597744 385026 597800
rect 385094 597744 385150 597800
rect 385218 597744 385274 597800
rect 385342 597744 385398 597800
rect 384970 586294 385026 586350
rect 385094 586294 385150 586350
rect 385218 586294 385274 586350
rect 385342 586294 385398 586350
rect 384970 586170 385026 586226
rect 385094 586170 385150 586226
rect 385218 586170 385274 586226
rect 385342 586170 385398 586226
rect 384970 586046 385026 586102
rect 385094 586046 385150 586102
rect 385218 586046 385274 586102
rect 385342 586046 385398 586102
rect 384970 585922 385026 585978
rect 385094 585922 385150 585978
rect 385218 585922 385274 585978
rect 385342 585922 385398 585978
rect 384970 568294 385026 568350
rect 385094 568294 385150 568350
rect 385218 568294 385274 568350
rect 385342 568294 385398 568350
rect 384970 568170 385026 568226
rect 385094 568170 385150 568226
rect 385218 568170 385274 568226
rect 385342 568170 385398 568226
rect 384970 568046 385026 568102
rect 385094 568046 385150 568102
rect 385218 568046 385274 568102
rect 385342 568046 385398 568102
rect 384970 567922 385026 567978
rect 385094 567922 385150 567978
rect 385218 567922 385274 567978
rect 385342 567922 385398 567978
rect 384970 550294 385026 550350
rect 385094 550294 385150 550350
rect 385218 550294 385274 550350
rect 385342 550294 385398 550350
rect 384970 550170 385026 550226
rect 385094 550170 385150 550226
rect 385218 550170 385274 550226
rect 385342 550170 385398 550226
rect 384970 550046 385026 550102
rect 385094 550046 385150 550102
rect 385218 550046 385274 550102
rect 385342 550046 385398 550102
rect 384970 549922 385026 549978
rect 385094 549922 385150 549978
rect 385218 549922 385274 549978
rect 385342 549922 385398 549978
rect 384970 532294 385026 532350
rect 385094 532294 385150 532350
rect 385218 532294 385274 532350
rect 385342 532294 385398 532350
rect 384970 532170 385026 532226
rect 385094 532170 385150 532226
rect 385218 532170 385274 532226
rect 385342 532170 385398 532226
rect 384970 532046 385026 532102
rect 385094 532046 385150 532102
rect 385218 532046 385274 532102
rect 385342 532046 385398 532102
rect 384970 531922 385026 531978
rect 385094 531922 385150 531978
rect 385218 531922 385274 531978
rect 385342 531922 385398 531978
rect 399250 597156 399306 597212
rect 399374 597156 399430 597212
rect 399498 597156 399554 597212
rect 399622 597156 399678 597212
rect 399250 597032 399306 597088
rect 399374 597032 399430 597088
rect 399498 597032 399554 597088
rect 399622 597032 399678 597088
rect 399250 596908 399306 596964
rect 399374 596908 399430 596964
rect 399498 596908 399554 596964
rect 399622 596908 399678 596964
rect 399250 596784 399306 596840
rect 399374 596784 399430 596840
rect 399498 596784 399554 596840
rect 399622 596784 399678 596840
rect 399250 580294 399306 580350
rect 399374 580294 399430 580350
rect 399498 580294 399554 580350
rect 399622 580294 399678 580350
rect 399250 580170 399306 580226
rect 399374 580170 399430 580226
rect 399498 580170 399554 580226
rect 399622 580170 399678 580226
rect 399250 580046 399306 580102
rect 399374 580046 399430 580102
rect 399498 580046 399554 580102
rect 399622 580046 399678 580102
rect 399250 579922 399306 579978
rect 399374 579922 399430 579978
rect 399498 579922 399554 579978
rect 399622 579922 399678 579978
rect 399250 562294 399306 562350
rect 399374 562294 399430 562350
rect 399498 562294 399554 562350
rect 399622 562294 399678 562350
rect 399250 562170 399306 562226
rect 399374 562170 399430 562226
rect 399498 562170 399554 562226
rect 399622 562170 399678 562226
rect 399250 562046 399306 562102
rect 399374 562046 399430 562102
rect 399498 562046 399554 562102
rect 399622 562046 399678 562102
rect 399250 561922 399306 561978
rect 399374 561922 399430 561978
rect 399498 561922 399554 561978
rect 399622 561922 399678 561978
rect 399250 544294 399306 544350
rect 399374 544294 399430 544350
rect 399498 544294 399554 544350
rect 399622 544294 399678 544350
rect 399250 544170 399306 544226
rect 399374 544170 399430 544226
rect 399498 544170 399554 544226
rect 399622 544170 399678 544226
rect 399250 544046 399306 544102
rect 399374 544046 399430 544102
rect 399498 544046 399554 544102
rect 399622 544046 399678 544102
rect 399250 543922 399306 543978
rect 399374 543922 399430 543978
rect 399498 543922 399554 543978
rect 399622 543922 399678 543978
rect 402970 598116 403026 598172
rect 403094 598116 403150 598172
rect 403218 598116 403274 598172
rect 403342 598116 403398 598172
rect 402970 597992 403026 598048
rect 403094 597992 403150 598048
rect 403218 597992 403274 598048
rect 403342 597992 403398 598048
rect 402970 597868 403026 597924
rect 403094 597868 403150 597924
rect 403218 597868 403274 597924
rect 403342 597868 403398 597924
rect 402970 597744 403026 597800
rect 403094 597744 403150 597800
rect 403218 597744 403274 597800
rect 403342 597744 403398 597800
rect 402970 586294 403026 586350
rect 403094 586294 403150 586350
rect 403218 586294 403274 586350
rect 403342 586294 403398 586350
rect 402970 586170 403026 586226
rect 403094 586170 403150 586226
rect 403218 586170 403274 586226
rect 403342 586170 403398 586226
rect 402970 586046 403026 586102
rect 403094 586046 403150 586102
rect 403218 586046 403274 586102
rect 403342 586046 403398 586102
rect 402970 585922 403026 585978
rect 403094 585922 403150 585978
rect 403218 585922 403274 585978
rect 403342 585922 403398 585978
rect 402970 568294 403026 568350
rect 403094 568294 403150 568350
rect 403218 568294 403274 568350
rect 403342 568294 403398 568350
rect 402970 568170 403026 568226
rect 403094 568170 403150 568226
rect 403218 568170 403274 568226
rect 403342 568170 403398 568226
rect 402970 568046 403026 568102
rect 403094 568046 403150 568102
rect 403218 568046 403274 568102
rect 403342 568046 403398 568102
rect 402970 567922 403026 567978
rect 403094 567922 403150 567978
rect 403218 567922 403274 567978
rect 403342 567922 403398 567978
rect 402970 550294 403026 550350
rect 403094 550294 403150 550350
rect 403218 550294 403274 550350
rect 403342 550294 403398 550350
rect 402970 550170 403026 550226
rect 403094 550170 403150 550226
rect 403218 550170 403274 550226
rect 403342 550170 403398 550226
rect 402970 550046 403026 550102
rect 403094 550046 403150 550102
rect 403218 550046 403274 550102
rect 403342 550046 403398 550102
rect 402970 549922 403026 549978
rect 403094 549922 403150 549978
rect 403218 549922 403274 549978
rect 403342 549922 403398 549978
rect 402970 532294 403026 532350
rect 403094 532294 403150 532350
rect 403218 532294 403274 532350
rect 403342 532294 403398 532350
rect 402970 532170 403026 532226
rect 403094 532170 403150 532226
rect 403218 532170 403274 532226
rect 403342 532170 403398 532226
rect 402970 532046 403026 532102
rect 403094 532046 403150 532102
rect 403218 532046 403274 532102
rect 403342 532046 403398 532102
rect 402970 531922 403026 531978
rect 403094 531922 403150 531978
rect 403218 531922 403274 531978
rect 403342 531922 403398 531978
rect 417250 597156 417306 597212
rect 417374 597156 417430 597212
rect 417498 597156 417554 597212
rect 417622 597156 417678 597212
rect 417250 597032 417306 597088
rect 417374 597032 417430 597088
rect 417498 597032 417554 597088
rect 417622 597032 417678 597088
rect 417250 596908 417306 596964
rect 417374 596908 417430 596964
rect 417498 596908 417554 596964
rect 417622 596908 417678 596964
rect 417250 596784 417306 596840
rect 417374 596784 417430 596840
rect 417498 596784 417554 596840
rect 417622 596784 417678 596840
rect 417250 580294 417306 580350
rect 417374 580294 417430 580350
rect 417498 580294 417554 580350
rect 417622 580294 417678 580350
rect 417250 580170 417306 580226
rect 417374 580170 417430 580226
rect 417498 580170 417554 580226
rect 417622 580170 417678 580226
rect 417250 580046 417306 580102
rect 417374 580046 417430 580102
rect 417498 580046 417554 580102
rect 417622 580046 417678 580102
rect 417250 579922 417306 579978
rect 417374 579922 417430 579978
rect 417498 579922 417554 579978
rect 417622 579922 417678 579978
rect 417250 562294 417306 562350
rect 417374 562294 417430 562350
rect 417498 562294 417554 562350
rect 417622 562294 417678 562350
rect 417250 562170 417306 562226
rect 417374 562170 417430 562226
rect 417498 562170 417554 562226
rect 417622 562170 417678 562226
rect 417250 562046 417306 562102
rect 417374 562046 417430 562102
rect 417498 562046 417554 562102
rect 417622 562046 417678 562102
rect 417250 561922 417306 561978
rect 417374 561922 417430 561978
rect 417498 561922 417554 561978
rect 417622 561922 417678 561978
rect 417250 544294 417306 544350
rect 417374 544294 417430 544350
rect 417498 544294 417554 544350
rect 417622 544294 417678 544350
rect 417250 544170 417306 544226
rect 417374 544170 417430 544226
rect 417498 544170 417554 544226
rect 417622 544170 417678 544226
rect 417250 544046 417306 544102
rect 417374 544046 417430 544102
rect 417498 544046 417554 544102
rect 417622 544046 417678 544102
rect 417250 543922 417306 543978
rect 417374 543922 417430 543978
rect 417498 543922 417554 543978
rect 417622 543922 417678 543978
rect 420970 598116 421026 598172
rect 421094 598116 421150 598172
rect 421218 598116 421274 598172
rect 421342 598116 421398 598172
rect 420970 597992 421026 598048
rect 421094 597992 421150 598048
rect 421218 597992 421274 598048
rect 421342 597992 421398 598048
rect 420970 597868 421026 597924
rect 421094 597868 421150 597924
rect 421218 597868 421274 597924
rect 421342 597868 421398 597924
rect 420970 597744 421026 597800
rect 421094 597744 421150 597800
rect 421218 597744 421274 597800
rect 421342 597744 421398 597800
rect 420970 586294 421026 586350
rect 421094 586294 421150 586350
rect 421218 586294 421274 586350
rect 421342 586294 421398 586350
rect 420970 586170 421026 586226
rect 421094 586170 421150 586226
rect 421218 586170 421274 586226
rect 421342 586170 421398 586226
rect 420970 586046 421026 586102
rect 421094 586046 421150 586102
rect 421218 586046 421274 586102
rect 421342 586046 421398 586102
rect 420970 585922 421026 585978
rect 421094 585922 421150 585978
rect 421218 585922 421274 585978
rect 421342 585922 421398 585978
rect 420970 568294 421026 568350
rect 421094 568294 421150 568350
rect 421218 568294 421274 568350
rect 421342 568294 421398 568350
rect 420970 568170 421026 568226
rect 421094 568170 421150 568226
rect 421218 568170 421274 568226
rect 421342 568170 421398 568226
rect 420970 568046 421026 568102
rect 421094 568046 421150 568102
rect 421218 568046 421274 568102
rect 421342 568046 421398 568102
rect 420970 567922 421026 567978
rect 421094 567922 421150 567978
rect 421218 567922 421274 567978
rect 421342 567922 421398 567978
rect 420970 550294 421026 550350
rect 421094 550294 421150 550350
rect 421218 550294 421274 550350
rect 421342 550294 421398 550350
rect 420970 550170 421026 550226
rect 421094 550170 421150 550226
rect 421218 550170 421274 550226
rect 421342 550170 421398 550226
rect 420970 550046 421026 550102
rect 421094 550046 421150 550102
rect 421218 550046 421274 550102
rect 421342 550046 421398 550102
rect 420970 549922 421026 549978
rect 421094 549922 421150 549978
rect 421218 549922 421274 549978
rect 421342 549922 421398 549978
rect 420970 532294 421026 532350
rect 421094 532294 421150 532350
rect 421218 532294 421274 532350
rect 421342 532294 421398 532350
rect 420970 532170 421026 532226
rect 421094 532170 421150 532226
rect 421218 532170 421274 532226
rect 421342 532170 421398 532226
rect 420970 532046 421026 532102
rect 421094 532046 421150 532102
rect 421218 532046 421274 532102
rect 421342 532046 421398 532102
rect 420970 531922 421026 531978
rect 421094 531922 421150 531978
rect 421218 531922 421274 531978
rect 421342 531922 421398 531978
rect 435250 597156 435306 597212
rect 435374 597156 435430 597212
rect 435498 597156 435554 597212
rect 435622 597156 435678 597212
rect 435250 597032 435306 597088
rect 435374 597032 435430 597088
rect 435498 597032 435554 597088
rect 435622 597032 435678 597088
rect 435250 596908 435306 596964
rect 435374 596908 435430 596964
rect 435498 596908 435554 596964
rect 435622 596908 435678 596964
rect 435250 596784 435306 596840
rect 435374 596784 435430 596840
rect 435498 596784 435554 596840
rect 435622 596784 435678 596840
rect 435250 580294 435306 580350
rect 435374 580294 435430 580350
rect 435498 580294 435554 580350
rect 435622 580294 435678 580350
rect 435250 580170 435306 580226
rect 435374 580170 435430 580226
rect 435498 580170 435554 580226
rect 435622 580170 435678 580226
rect 435250 580046 435306 580102
rect 435374 580046 435430 580102
rect 435498 580046 435554 580102
rect 435622 580046 435678 580102
rect 435250 579922 435306 579978
rect 435374 579922 435430 579978
rect 435498 579922 435554 579978
rect 435622 579922 435678 579978
rect 435250 562294 435306 562350
rect 435374 562294 435430 562350
rect 435498 562294 435554 562350
rect 435622 562294 435678 562350
rect 435250 562170 435306 562226
rect 435374 562170 435430 562226
rect 435498 562170 435554 562226
rect 435622 562170 435678 562226
rect 435250 562046 435306 562102
rect 435374 562046 435430 562102
rect 435498 562046 435554 562102
rect 435622 562046 435678 562102
rect 435250 561922 435306 561978
rect 435374 561922 435430 561978
rect 435498 561922 435554 561978
rect 435622 561922 435678 561978
rect 435250 544294 435306 544350
rect 435374 544294 435430 544350
rect 435498 544294 435554 544350
rect 435622 544294 435678 544350
rect 435250 544170 435306 544226
rect 435374 544170 435430 544226
rect 435498 544170 435554 544226
rect 435622 544170 435678 544226
rect 435250 544046 435306 544102
rect 435374 544046 435430 544102
rect 435498 544046 435554 544102
rect 435622 544046 435678 544102
rect 435250 543922 435306 543978
rect 435374 543922 435430 543978
rect 435498 543922 435554 543978
rect 435622 543922 435678 543978
rect 438970 598116 439026 598172
rect 439094 598116 439150 598172
rect 439218 598116 439274 598172
rect 439342 598116 439398 598172
rect 438970 597992 439026 598048
rect 439094 597992 439150 598048
rect 439218 597992 439274 598048
rect 439342 597992 439398 598048
rect 438970 597868 439026 597924
rect 439094 597868 439150 597924
rect 439218 597868 439274 597924
rect 439342 597868 439398 597924
rect 438970 597744 439026 597800
rect 439094 597744 439150 597800
rect 439218 597744 439274 597800
rect 439342 597744 439398 597800
rect 438970 586294 439026 586350
rect 439094 586294 439150 586350
rect 439218 586294 439274 586350
rect 439342 586294 439398 586350
rect 438970 586170 439026 586226
rect 439094 586170 439150 586226
rect 439218 586170 439274 586226
rect 439342 586170 439398 586226
rect 438970 586046 439026 586102
rect 439094 586046 439150 586102
rect 439218 586046 439274 586102
rect 439342 586046 439398 586102
rect 438970 585922 439026 585978
rect 439094 585922 439150 585978
rect 439218 585922 439274 585978
rect 439342 585922 439398 585978
rect 438970 568294 439026 568350
rect 439094 568294 439150 568350
rect 439218 568294 439274 568350
rect 439342 568294 439398 568350
rect 438970 568170 439026 568226
rect 439094 568170 439150 568226
rect 439218 568170 439274 568226
rect 439342 568170 439398 568226
rect 438970 568046 439026 568102
rect 439094 568046 439150 568102
rect 439218 568046 439274 568102
rect 439342 568046 439398 568102
rect 438970 567922 439026 567978
rect 439094 567922 439150 567978
rect 439218 567922 439274 567978
rect 439342 567922 439398 567978
rect 438970 550294 439026 550350
rect 439094 550294 439150 550350
rect 439218 550294 439274 550350
rect 439342 550294 439398 550350
rect 438970 550170 439026 550226
rect 439094 550170 439150 550226
rect 439218 550170 439274 550226
rect 439342 550170 439398 550226
rect 438970 550046 439026 550102
rect 439094 550046 439150 550102
rect 439218 550046 439274 550102
rect 439342 550046 439398 550102
rect 438970 549922 439026 549978
rect 439094 549922 439150 549978
rect 439218 549922 439274 549978
rect 439342 549922 439398 549978
rect 438970 532294 439026 532350
rect 439094 532294 439150 532350
rect 439218 532294 439274 532350
rect 439342 532294 439398 532350
rect 438970 532170 439026 532226
rect 439094 532170 439150 532226
rect 439218 532170 439274 532226
rect 439342 532170 439398 532226
rect 438970 532046 439026 532102
rect 439094 532046 439150 532102
rect 439218 532046 439274 532102
rect 439342 532046 439398 532102
rect 438970 531922 439026 531978
rect 439094 531922 439150 531978
rect 439218 531922 439274 531978
rect 439342 531922 439398 531978
rect 453250 597156 453306 597212
rect 453374 597156 453430 597212
rect 453498 597156 453554 597212
rect 453622 597156 453678 597212
rect 453250 597032 453306 597088
rect 453374 597032 453430 597088
rect 453498 597032 453554 597088
rect 453622 597032 453678 597088
rect 453250 596908 453306 596964
rect 453374 596908 453430 596964
rect 453498 596908 453554 596964
rect 453622 596908 453678 596964
rect 453250 596784 453306 596840
rect 453374 596784 453430 596840
rect 453498 596784 453554 596840
rect 453622 596784 453678 596840
rect 453250 580294 453306 580350
rect 453374 580294 453430 580350
rect 453498 580294 453554 580350
rect 453622 580294 453678 580350
rect 453250 580170 453306 580226
rect 453374 580170 453430 580226
rect 453498 580170 453554 580226
rect 453622 580170 453678 580226
rect 453250 580046 453306 580102
rect 453374 580046 453430 580102
rect 453498 580046 453554 580102
rect 453622 580046 453678 580102
rect 453250 579922 453306 579978
rect 453374 579922 453430 579978
rect 453498 579922 453554 579978
rect 453622 579922 453678 579978
rect 453250 562294 453306 562350
rect 453374 562294 453430 562350
rect 453498 562294 453554 562350
rect 453622 562294 453678 562350
rect 453250 562170 453306 562226
rect 453374 562170 453430 562226
rect 453498 562170 453554 562226
rect 453622 562170 453678 562226
rect 453250 562046 453306 562102
rect 453374 562046 453430 562102
rect 453498 562046 453554 562102
rect 453622 562046 453678 562102
rect 453250 561922 453306 561978
rect 453374 561922 453430 561978
rect 453498 561922 453554 561978
rect 453622 561922 453678 561978
rect 453250 544294 453306 544350
rect 453374 544294 453430 544350
rect 453498 544294 453554 544350
rect 453622 544294 453678 544350
rect 453250 544170 453306 544226
rect 453374 544170 453430 544226
rect 453498 544170 453554 544226
rect 453622 544170 453678 544226
rect 453250 544046 453306 544102
rect 453374 544046 453430 544102
rect 453498 544046 453554 544102
rect 453622 544046 453678 544102
rect 453250 543922 453306 543978
rect 453374 543922 453430 543978
rect 453498 543922 453554 543978
rect 453622 543922 453678 543978
rect 456970 598116 457026 598172
rect 457094 598116 457150 598172
rect 457218 598116 457274 598172
rect 457342 598116 457398 598172
rect 456970 597992 457026 598048
rect 457094 597992 457150 598048
rect 457218 597992 457274 598048
rect 457342 597992 457398 598048
rect 456970 597868 457026 597924
rect 457094 597868 457150 597924
rect 457218 597868 457274 597924
rect 457342 597868 457398 597924
rect 456970 597744 457026 597800
rect 457094 597744 457150 597800
rect 457218 597744 457274 597800
rect 457342 597744 457398 597800
rect 456970 586294 457026 586350
rect 457094 586294 457150 586350
rect 457218 586294 457274 586350
rect 457342 586294 457398 586350
rect 456970 586170 457026 586226
rect 457094 586170 457150 586226
rect 457218 586170 457274 586226
rect 457342 586170 457398 586226
rect 456970 586046 457026 586102
rect 457094 586046 457150 586102
rect 457218 586046 457274 586102
rect 457342 586046 457398 586102
rect 456970 585922 457026 585978
rect 457094 585922 457150 585978
rect 457218 585922 457274 585978
rect 457342 585922 457398 585978
rect 456970 568294 457026 568350
rect 457094 568294 457150 568350
rect 457218 568294 457274 568350
rect 457342 568294 457398 568350
rect 456970 568170 457026 568226
rect 457094 568170 457150 568226
rect 457218 568170 457274 568226
rect 457342 568170 457398 568226
rect 456970 568046 457026 568102
rect 457094 568046 457150 568102
rect 457218 568046 457274 568102
rect 457342 568046 457398 568102
rect 456970 567922 457026 567978
rect 457094 567922 457150 567978
rect 457218 567922 457274 567978
rect 457342 567922 457398 567978
rect 456970 550294 457026 550350
rect 457094 550294 457150 550350
rect 457218 550294 457274 550350
rect 457342 550294 457398 550350
rect 456970 550170 457026 550226
rect 457094 550170 457150 550226
rect 457218 550170 457274 550226
rect 457342 550170 457398 550226
rect 456970 550046 457026 550102
rect 457094 550046 457150 550102
rect 457218 550046 457274 550102
rect 457342 550046 457398 550102
rect 456970 549922 457026 549978
rect 457094 549922 457150 549978
rect 457218 549922 457274 549978
rect 457342 549922 457398 549978
rect 456970 532294 457026 532350
rect 457094 532294 457150 532350
rect 457218 532294 457274 532350
rect 457342 532294 457398 532350
rect 456970 532170 457026 532226
rect 457094 532170 457150 532226
rect 457218 532170 457274 532226
rect 457342 532170 457398 532226
rect 456970 532046 457026 532102
rect 457094 532046 457150 532102
rect 457218 532046 457274 532102
rect 457342 532046 457398 532102
rect 456970 531922 457026 531978
rect 457094 531922 457150 531978
rect 457218 531922 457274 531978
rect 457342 531922 457398 531978
rect 471250 597156 471306 597212
rect 471374 597156 471430 597212
rect 471498 597156 471554 597212
rect 471622 597156 471678 597212
rect 471250 597032 471306 597088
rect 471374 597032 471430 597088
rect 471498 597032 471554 597088
rect 471622 597032 471678 597088
rect 471250 596908 471306 596964
rect 471374 596908 471430 596964
rect 471498 596908 471554 596964
rect 471622 596908 471678 596964
rect 471250 596784 471306 596840
rect 471374 596784 471430 596840
rect 471498 596784 471554 596840
rect 471622 596784 471678 596840
rect 471250 580294 471306 580350
rect 471374 580294 471430 580350
rect 471498 580294 471554 580350
rect 471622 580294 471678 580350
rect 471250 580170 471306 580226
rect 471374 580170 471430 580226
rect 471498 580170 471554 580226
rect 471622 580170 471678 580226
rect 471250 580046 471306 580102
rect 471374 580046 471430 580102
rect 471498 580046 471554 580102
rect 471622 580046 471678 580102
rect 471250 579922 471306 579978
rect 471374 579922 471430 579978
rect 471498 579922 471554 579978
rect 471622 579922 471678 579978
rect 471250 562294 471306 562350
rect 471374 562294 471430 562350
rect 471498 562294 471554 562350
rect 471622 562294 471678 562350
rect 471250 562170 471306 562226
rect 471374 562170 471430 562226
rect 471498 562170 471554 562226
rect 471622 562170 471678 562226
rect 471250 562046 471306 562102
rect 471374 562046 471430 562102
rect 471498 562046 471554 562102
rect 471622 562046 471678 562102
rect 471250 561922 471306 561978
rect 471374 561922 471430 561978
rect 471498 561922 471554 561978
rect 471622 561922 471678 561978
rect 471250 544294 471306 544350
rect 471374 544294 471430 544350
rect 471498 544294 471554 544350
rect 471622 544294 471678 544350
rect 471250 544170 471306 544226
rect 471374 544170 471430 544226
rect 471498 544170 471554 544226
rect 471622 544170 471678 544226
rect 471250 544046 471306 544102
rect 471374 544046 471430 544102
rect 471498 544046 471554 544102
rect 471622 544046 471678 544102
rect 471250 543922 471306 543978
rect 471374 543922 471430 543978
rect 471498 543922 471554 543978
rect 471622 543922 471678 543978
rect 474970 598116 475026 598172
rect 475094 598116 475150 598172
rect 475218 598116 475274 598172
rect 475342 598116 475398 598172
rect 474970 597992 475026 598048
rect 475094 597992 475150 598048
rect 475218 597992 475274 598048
rect 475342 597992 475398 598048
rect 474970 597868 475026 597924
rect 475094 597868 475150 597924
rect 475218 597868 475274 597924
rect 475342 597868 475398 597924
rect 474970 597744 475026 597800
rect 475094 597744 475150 597800
rect 475218 597744 475274 597800
rect 475342 597744 475398 597800
rect 474970 586294 475026 586350
rect 475094 586294 475150 586350
rect 475218 586294 475274 586350
rect 475342 586294 475398 586350
rect 474970 586170 475026 586226
rect 475094 586170 475150 586226
rect 475218 586170 475274 586226
rect 475342 586170 475398 586226
rect 474970 586046 475026 586102
rect 475094 586046 475150 586102
rect 475218 586046 475274 586102
rect 475342 586046 475398 586102
rect 474970 585922 475026 585978
rect 475094 585922 475150 585978
rect 475218 585922 475274 585978
rect 475342 585922 475398 585978
rect 474970 568294 475026 568350
rect 475094 568294 475150 568350
rect 475218 568294 475274 568350
rect 475342 568294 475398 568350
rect 474970 568170 475026 568226
rect 475094 568170 475150 568226
rect 475218 568170 475274 568226
rect 475342 568170 475398 568226
rect 474970 568046 475026 568102
rect 475094 568046 475150 568102
rect 475218 568046 475274 568102
rect 475342 568046 475398 568102
rect 474970 567922 475026 567978
rect 475094 567922 475150 567978
rect 475218 567922 475274 567978
rect 475342 567922 475398 567978
rect 474970 550294 475026 550350
rect 475094 550294 475150 550350
rect 475218 550294 475274 550350
rect 475342 550294 475398 550350
rect 474970 550170 475026 550226
rect 475094 550170 475150 550226
rect 475218 550170 475274 550226
rect 475342 550170 475398 550226
rect 474970 550046 475026 550102
rect 475094 550046 475150 550102
rect 475218 550046 475274 550102
rect 475342 550046 475398 550102
rect 474970 549922 475026 549978
rect 475094 549922 475150 549978
rect 475218 549922 475274 549978
rect 475342 549922 475398 549978
rect 474970 532294 475026 532350
rect 475094 532294 475150 532350
rect 475218 532294 475274 532350
rect 475342 532294 475398 532350
rect 474970 532170 475026 532226
rect 475094 532170 475150 532226
rect 475218 532170 475274 532226
rect 475342 532170 475398 532226
rect 474970 532046 475026 532102
rect 475094 532046 475150 532102
rect 475218 532046 475274 532102
rect 475342 532046 475398 532102
rect 474970 531922 475026 531978
rect 475094 531922 475150 531978
rect 475218 531922 475274 531978
rect 475342 531922 475398 531978
rect 489250 597156 489306 597212
rect 489374 597156 489430 597212
rect 489498 597156 489554 597212
rect 489622 597156 489678 597212
rect 489250 597032 489306 597088
rect 489374 597032 489430 597088
rect 489498 597032 489554 597088
rect 489622 597032 489678 597088
rect 489250 596908 489306 596964
rect 489374 596908 489430 596964
rect 489498 596908 489554 596964
rect 489622 596908 489678 596964
rect 489250 596784 489306 596840
rect 489374 596784 489430 596840
rect 489498 596784 489554 596840
rect 489622 596784 489678 596840
rect 489250 580294 489306 580350
rect 489374 580294 489430 580350
rect 489498 580294 489554 580350
rect 489622 580294 489678 580350
rect 489250 580170 489306 580226
rect 489374 580170 489430 580226
rect 489498 580170 489554 580226
rect 489622 580170 489678 580226
rect 489250 580046 489306 580102
rect 489374 580046 489430 580102
rect 489498 580046 489554 580102
rect 489622 580046 489678 580102
rect 489250 579922 489306 579978
rect 489374 579922 489430 579978
rect 489498 579922 489554 579978
rect 489622 579922 489678 579978
rect 489250 562294 489306 562350
rect 489374 562294 489430 562350
rect 489498 562294 489554 562350
rect 489622 562294 489678 562350
rect 489250 562170 489306 562226
rect 489374 562170 489430 562226
rect 489498 562170 489554 562226
rect 489622 562170 489678 562226
rect 489250 562046 489306 562102
rect 489374 562046 489430 562102
rect 489498 562046 489554 562102
rect 489622 562046 489678 562102
rect 489250 561922 489306 561978
rect 489374 561922 489430 561978
rect 489498 561922 489554 561978
rect 489622 561922 489678 561978
rect 489250 544294 489306 544350
rect 489374 544294 489430 544350
rect 489498 544294 489554 544350
rect 489622 544294 489678 544350
rect 489250 544170 489306 544226
rect 489374 544170 489430 544226
rect 489498 544170 489554 544226
rect 489622 544170 489678 544226
rect 489250 544046 489306 544102
rect 489374 544046 489430 544102
rect 489498 544046 489554 544102
rect 489622 544046 489678 544102
rect 489250 543922 489306 543978
rect 489374 543922 489430 543978
rect 489498 543922 489554 543978
rect 489622 543922 489678 543978
rect 492970 598116 493026 598172
rect 493094 598116 493150 598172
rect 493218 598116 493274 598172
rect 493342 598116 493398 598172
rect 492970 597992 493026 598048
rect 493094 597992 493150 598048
rect 493218 597992 493274 598048
rect 493342 597992 493398 598048
rect 492970 597868 493026 597924
rect 493094 597868 493150 597924
rect 493218 597868 493274 597924
rect 493342 597868 493398 597924
rect 492970 597744 493026 597800
rect 493094 597744 493150 597800
rect 493218 597744 493274 597800
rect 493342 597744 493398 597800
rect 492970 586294 493026 586350
rect 493094 586294 493150 586350
rect 493218 586294 493274 586350
rect 493342 586294 493398 586350
rect 492970 586170 493026 586226
rect 493094 586170 493150 586226
rect 493218 586170 493274 586226
rect 493342 586170 493398 586226
rect 492970 586046 493026 586102
rect 493094 586046 493150 586102
rect 493218 586046 493274 586102
rect 493342 586046 493398 586102
rect 492970 585922 493026 585978
rect 493094 585922 493150 585978
rect 493218 585922 493274 585978
rect 493342 585922 493398 585978
rect 492970 568294 493026 568350
rect 493094 568294 493150 568350
rect 493218 568294 493274 568350
rect 493342 568294 493398 568350
rect 492970 568170 493026 568226
rect 493094 568170 493150 568226
rect 493218 568170 493274 568226
rect 493342 568170 493398 568226
rect 492970 568046 493026 568102
rect 493094 568046 493150 568102
rect 493218 568046 493274 568102
rect 493342 568046 493398 568102
rect 492970 567922 493026 567978
rect 493094 567922 493150 567978
rect 493218 567922 493274 567978
rect 493342 567922 493398 567978
rect 492970 550294 493026 550350
rect 493094 550294 493150 550350
rect 493218 550294 493274 550350
rect 493342 550294 493398 550350
rect 492970 550170 493026 550226
rect 493094 550170 493150 550226
rect 493218 550170 493274 550226
rect 493342 550170 493398 550226
rect 492970 550046 493026 550102
rect 493094 550046 493150 550102
rect 493218 550046 493274 550102
rect 493342 550046 493398 550102
rect 492970 549922 493026 549978
rect 493094 549922 493150 549978
rect 493218 549922 493274 549978
rect 493342 549922 493398 549978
rect 492970 532294 493026 532350
rect 493094 532294 493150 532350
rect 493218 532294 493274 532350
rect 493342 532294 493398 532350
rect 492970 532170 493026 532226
rect 493094 532170 493150 532226
rect 493218 532170 493274 532226
rect 493342 532170 493398 532226
rect 492970 532046 493026 532102
rect 493094 532046 493150 532102
rect 493218 532046 493274 532102
rect 493342 532046 493398 532102
rect 492970 531922 493026 531978
rect 493094 531922 493150 531978
rect 493218 531922 493274 531978
rect 493342 531922 493398 531978
rect 507250 597156 507306 597212
rect 507374 597156 507430 597212
rect 507498 597156 507554 597212
rect 507622 597156 507678 597212
rect 507250 597032 507306 597088
rect 507374 597032 507430 597088
rect 507498 597032 507554 597088
rect 507622 597032 507678 597088
rect 507250 596908 507306 596964
rect 507374 596908 507430 596964
rect 507498 596908 507554 596964
rect 507622 596908 507678 596964
rect 507250 596784 507306 596840
rect 507374 596784 507430 596840
rect 507498 596784 507554 596840
rect 507622 596784 507678 596840
rect 507250 580294 507306 580350
rect 507374 580294 507430 580350
rect 507498 580294 507554 580350
rect 507622 580294 507678 580350
rect 507250 580170 507306 580226
rect 507374 580170 507430 580226
rect 507498 580170 507554 580226
rect 507622 580170 507678 580226
rect 507250 580046 507306 580102
rect 507374 580046 507430 580102
rect 507498 580046 507554 580102
rect 507622 580046 507678 580102
rect 507250 579922 507306 579978
rect 507374 579922 507430 579978
rect 507498 579922 507554 579978
rect 507622 579922 507678 579978
rect 507250 562294 507306 562350
rect 507374 562294 507430 562350
rect 507498 562294 507554 562350
rect 507622 562294 507678 562350
rect 507250 562170 507306 562226
rect 507374 562170 507430 562226
rect 507498 562170 507554 562226
rect 507622 562170 507678 562226
rect 507250 562046 507306 562102
rect 507374 562046 507430 562102
rect 507498 562046 507554 562102
rect 507622 562046 507678 562102
rect 507250 561922 507306 561978
rect 507374 561922 507430 561978
rect 507498 561922 507554 561978
rect 507622 561922 507678 561978
rect 507250 544294 507306 544350
rect 507374 544294 507430 544350
rect 507498 544294 507554 544350
rect 507622 544294 507678 544350
rect 507250 544170 507306 544226
rect 507374 544170 507430 544226
rect 507498 544170 507554 544226
rect 507622 544170 507678 544226
rect 507250 544046 507306 544102
rect 507374 544046 507430 544102
rect 507498 544046 507554 544102
rect 507622 544046 507678 544102
rect 507250 543922 507306 543978
rect 507374 543922 507430 543978
rect 507498 543922 507554 543978
rect 507622 543922 507678 543978
rect 510970 598116 511026 598172
rect 511094 598116 511150 598172
rect 511218 598116 511274 598172
rect 511342 598116 511398 598172
rect 510970 597992 511026 598048
rect 511094 597992 511150 598048
rect 511218 597992 511274 598048
rect 511342 597992 511398 598048
rect 510970 597868 511026 597924
rect 511094 597868 511150 597924
rect 511218 597868 511274 597924
rect 511342 597868 511398 597924
rect 510970 597744 511026 597800
rect 511094 597744 511150 597800
rect 511218 597744 511274 597800
rect 511342 597744 511398 597800
rect 510970 586294 511026 586350
rect 511094 586294 511150 586350
rect 511218 586294 511274 586350
rect 511342 586294 511398 586350
rect 510970 586170 511026 586226
rect 511094 586170 511150 586226
rect 511218 586170 511274 586226
rect 511342 586170 511398 586226
rect 510970 586046 511026 586102
rect 511094 586046 511150 586102
rect 511218 586046 511274 586102
rect 511342 586046 511398 586102
rect 510970 585922 511026 585978
rect 511094 585922 511150 585978
rect 511218 585922 511274 585978
rect 511342 585922 511398 585978
rect 510970 568294 511026 568350
rect 511094 568294 511150 568350
rect 511218 568294 511274 568350
rect 511342 568294 511398 568350
rect 510970 568170 511026 568226
rect 511094 568170 511150 568226
rect 511218 568170 511274 568226
rect 511342 568170 511398 568226
rect 510970 568046 511026 568102
rect 511094 568046 511150 568102
rect 511218 568046 511274 568102
rect 511342 568046 511398 568102
rect 510970 567922 511026 567978
rect 511094 567922 511150 567978
rect 511218 567922 511274 567978
rect 511342 567922 511398 567978
rect 510970 550294 511026 550350
rect 511094 550294 511150 550350
rect 511218 550294 511274 550350
rect 511342 550294 511398 550350
rect 510970 550170 511026 550226
rect 511094 550170 511150 550226
rect 511218 550170 511274 550226
rect 511342 550170 511398 550226
rect 510970 550046 511026 550102
rect 511094 550046 511150 550102
rect 511218 550046 511274 550102
rect 511342 550046 511398 550102
rect 510970 549922 511026 549978
rect 511094 549922 511150 549978
rect 511218 549922 511274 549978
rect 511342 549922 511398 549978
rect 510970 532294 511026 532350
rect 511094 532294 511150 532350
rect 511218 532294 511274 532350
rect 511342 532294 511398 532350
rect 510970 532170 511026 532226
rect 511094 532170 511150 532226
rect 511218 532170 511274 532226
rect 511342 532170 511398 532226
rect 510970 532046 511026 532102
rect 511094 532046 511150 532102
rect 511218 532046 511274 532102
rect 511342 532046 511398 532102
rect 510970 531922 511026 531978
rect 511094 531922 511150 531978
rect 511218 531922 511274 531978
rect 511342 531922 511398 531978
rect 525250 597156 525306 597212
rect 525374 597156 525430 597212
rect 525498 597156 525554 597212
rect 525622 597156 525678 597212
rect 525250 597032 525306 597088
rect 525374 597032 525430 597088
rect 525498 597032 525554 597088
rect 525622 597032 525678 597088
rect 525250 596908 525306 596964
rect 525374 596908 525430 596964
rect 525498 596908 525554 596964
rect 525622 596908 525678 596964
rect 525250 596784 525306 596840
rect 525374 596784 525430 596840
rect 525498 596784 525554 596840
rect 525622 596784 525678 596840
rect 525250 580294 525306 580350
rect 525374 580294 525430 580350
rect 525498 580294 525554 580350
rect 525622 580294 525678 580350
rect 525250 580170 525306 580226
rect 525374 580170 525430 580226
rect 525498 580170 525554 580226
rect 525622 580170 525678 580226
rect 525250 580046 525306 580102
rect 525374 580046 525430 580102
rect 525498 580046 525554 580102
rect 525622 580046 525678 580102
rect 525250 579922 525306 579978
rect 525374 579922 525430 579978
rect 525498 579922 525554 579978
rect 525622 579922 525678 579978
rect 525250 562294 525306 562350
rect 525374 562294 525430 562350
rect 525498 562294 525554 562350
rect 525622 562294 525678 562350
rect 525250 562170 525306 562226
rect 525374 562170 525430 562226
rect 525498 562170 525554 562226
rect 525622 562170 525678 562226
rect 525250 562046 525306 562102
rect 525374 562046 525430 562102
rect 525498 562046 525554 562102
rect 525622 562046 525678 562102
rect 525250 561922 525306 561978
rect 525374 561922 525430 561978
rect 525498 561922 525554 561978
rect 525622 561922 525678 561978
rect 525250 544294 525306 544350
rect 525374 544294 525430 544350
rect 525498 544294 525554 544350
rect 525622 544294 525678 544350
rect 525250 544170 525306 544226
rect 525374 544170 525430 544226
rect 525498 544170 525554 544226
rect 525622 544170 525678 544226
rect 525250 544046 525306 544102
rect 525374 544046 525430 544102
rect 525498 544046 525554 544102
rect 525622 544046 525678 544102
rect 525250 543922 525306 543978
rect 525374 543922 525430 543978
rect 525498 543922 525554 543978
rect 525622 543922 525678 543978
rect 528970 598116 529026 598172
rect 529094 598116 529150 598172
rect 529218 598116 529274 598172
rect 529342 598116 529398 598172
rect 528970 597992 529026 598048
rect 529094 597992 529150 598048
rect 529218 597992 529274 598048
rect 529342 597992 529398 598048
rect 528970 597868 529026 597924
rect 529094 597868 529150 597924
rect 529218 597868 529274 597924
rect 529342 597868 529398 597924
rect 528970 597744 529026 597800
rect 529094 597744 529150 597800
rect 529218 597744 529274 597800
rect 529342 597744 529398 597800
rect 528970 586294 529026 586350
rect 529094 586294 529150 586350
rect 529218 586294 529274 586350
rect 529342 586294 529398 586350
rect 528970 586170 529026 586226
rect 529094 586170 529150 586226
rect 529218 586170 529274 586226
rect 529342 586170 529398 586226
rect 528970 586046 529026 586102
rect 529094 586046 529150 586102
rect 529218 586046 529274 586102
rect 529342 586046 529398 586102
rect 528970 585922 529026 585978
rect 529094 585922 529150 585978
rect 529218 585922 529274 585978
rect 529342 585922 529398 585978
rect 528970 568294 529026 568350
rect 529094 568294 529150 568350
rect 529218 568294 529274 568350
rect 529342 568294 529398 568350
rect 528970 568170 529026 568226
rect 529094 568170 529150 568226
rect 529218 568170 529274 568226
rect 529342 568170 529398 568226
rect 528970 568046 529026 568102
rect 529094 568046 529150 568102
rect 529218 568046 529274 568102
rect 529342 568046 529398 568102
rect 528970 567922 529026 567978
rect 529094 567922 529150 567978
rect 529218 567922 529274 567978
rect 529342 567922 529398 567978
rect 528970 550294 529026 550350
rect 529094 550294 529150 550350
rect 529218 550294 529274 550350
rect 529342 550294 529398 550350
rect 528970 550170 529026 550226
rect 529094 550170 529150 550226
rect 529218 550170 529274 550226
rect 529342 550170 529398 550226
rect 528970 550046 529026 550102
rect 529094 550046 529150 550102
rect 529218 550046 529274 550102
rect 529342 550046 529398 550102
rect 528970 549922 529026 549978
rect 529094 549922 529150 549978
rect 529218 549922 529274 549978
rect 529342 549922 529398 549978
rect 528970 532294 529026 532350
rect 529094 532294 529150 532350
rect 529218 532294 529274 532350
rect 529342 532294 529398 532350
rect 528970 532170 529026 532226
rect 529094 532170 529150 532226
rect 529218 532170 529274 532226
rect 529342 532170 529398 532226
rect 528970 532046 529026 532102
rect 529094 532046 529150 532102
rect 529218 532046 529274 532102
rect 529342 532046 529398 532102
rect 528970 531922 529026 531978
rect 529094 531922 529150 531978
rect 529218 531922 529274 531978
rect 529342 531922 529398 531978
rect 543250 597156 543306 597212
rect 543374 597156 543430 597212
rect 543498 597156 543554 597212
rect 543622 597156 543678 597212
rect 543250 597032 543306 597088
rect 543374 597032 543430 597088
rect 543498 597032 543554 597088
rect 543622 597032 543678 597088
rect 543250 596908 543306 596964
rect 543374 596908 543430 596964
rect 543498 596908 543554 596964
rect 543622 596908 543678 596964
rect 543250 596784 543306 596840
rect 543374 596784 543430 596840
rect 543498 596784 543554 596840
rect 543622 596784 543678 596840
rect 543250 580294 543306 580350
rect 543374 580294 543430 580350
rect 543498 580294 543554 580350
rect 543622 580294 543678 580350
rect 543250 580170 543306 580226
rect 543374 580170 543430 580226
rect 543498 580170 543554 580226
rect 543622 580170 543678 580226
rect 543250 580046 543306 580102
rect 543374 580046 543430 580102
rect 543498 580046 543554 580102
rect 543622 580046 543678 580102
rect 543250 579922 543306 579978
rect 543374 579922 543430 579978
rect 543498 579922 543554 579978
rect 543622 579922 543678 579978
rect 543250 562294 543306 562350
rect 543374 562294 543430 562350
rect 543498 562294 543554 562350
rect 543622 562294 543678 562350
rect 543250 562170 543306 562226
rect 543374 562170 543430 562226
rect 543498 562170 543554 562226
rect 543622 562170 543678 562226
rect 543250 562046 543306 562102
rect 543374 562046 543430 562102
rect 543498 562046 543554 562102
rect 543622 562046 543678 562102
rect 543250 561922 543306 561978
rect 543374 561922 543430 561978
rect 543498 561922 543554 561978
rect 543622 561922 543678 561978
rect 543250 544294 543306 544350
rect 543374 544294 543430 544350
rect 543498 544294 543554 544350
rect 543622 544294 543678 544350
rect 543250 544170 543306 544226
rect 543374 544170 543430 544226
rect 543498 544170 543554 544226
rect 543622 544170 543678 544226
rect 543250 544046 543306 544102
rect 543374 544046 543430 544102
rect 543498 544046 543554 544102
rect 543622 544046 543678 544102
rect 543250 543922 543306 543978
rect 543374 543922 543430 543978
rect 543498 543922 543554 543978
rect 543622 543922 543678 543978
rect 546970 598116 547026 598172
rect 547094 598116 547150 598172
rect 547218 598116 547274 598172
rect 547342 598116 547398 598172
rect 546970 597992 547026 598048
rect 547094 597992 547150 598048
rect 547218 597992 547274 598048
rect 547342 597992 547398 598048
rect 546970 597868 547026 597924
rect 547094 597868 547150 597924
rect 547218 597868 547274 597924
rect 547342 597868 547398 597924
rect 546970 597744 547026 597800
rect 547094 597744 547150 597800
rect 547218 597744 547274 597800
rect 547342 597744 547398 597800
rect 546970 586294 547026 586350
rect 547094 586294 547150 586350
rect 547218 586294 547274 586350
rect 547342 586294 547398 586350
rect 546970 586170 547026 586226
rect 547094 586170 547150 586226
rect 547218 586170 547274 586226
rect 547342 586170 547398 586226
rect 546970 586046 547026 586102
rect 547094 586046 547150 586102
rect 547218 586046 547274 586102
rect 547342 586046 547398 586102
rect 546970 585922 547026 585978
rect 547094 585922 547150 585978
rect 547218 585922 547274 585978
rect 547342 585922 547398 585978
rect 546970 568294 547026 568350
rect 547094 568294 547150 568350
rect 547218 568294 547274 568350
rect 547342 568294 547398 568350
rect 546970 568170 547026 568226
rect 547094 568170 547150 568226
rect 547218 568170 547274 568226
rect 547342 568170 547398 568226
rect 546970 568046 547026 568102
rect 547094 568046 547150 568102
rect 547218 568046 547274 568102
rect 547342 568046 547398 568102
rect 546970 567922 547026 567978
rect 547094 567922 547150 567978
rect 547218 567922 547274 567978
rect 547342 567922 547398 567978
rect 546970 550294 547026 550350
rect 547094 550294 547150 550350
rect 547218 550294 547274 550350
rect 547342 550294 547398 550350
rect 546970 550170 547026 550226
rect 547094 550170 547150 550226
rect 547218 550170 547274 550226
rect 547342 550170 547398 550226
rect 546970 550046 547026 550102
rect 547094 550046 547150 550102
rect 547218 550046 547274 550102
rect 547342 550046 547398 550102
rect 546970 549922 547026 549978
rect 547094 549922 547150 549978
rect 547218 549922 547274 549978
rect 547342 549922 547398 549978
rect 546970 532294 547026 532350
rect 547094 532294 547150 532350
rect 547218 532294 547274 532350
rect 547342 532294 547398 532350
rect 546970 532170 547026 532226
rect 547094 532170 547150 532226
rect 547218 532170 547274 532226
rect 547342 532170 547398 532226
rect 546970 532046 547026 532102
rect 547094 532046 547150 532102
rect 547218 532046 547274 532102
rect 547342 532046 547398 532102
rect 546970 531922 547026 531978
rect 547094 531922 547150 531978
rect 547218 531922 547274 531978
rect 547342 531922 547398 531978
rect 561250 597156 561306 597212
rect 561374 597156 561430 597212
rect 561498 597156 561554 597212
rect 561622 597156 561678 597212
rect 561250 597032 561306 597088
rect 561374 597032 561430 597088
rect 561498 597032 561554 597088
rect 561622 597032 561678 597088
rect 561250 596908 561306 596964
rect 561374 596908 561430 596964
rect 561498 596908 561554 596964
rect 561622 596908 561678 596964
rect 561250 596784 561306 596840
rect 561374 596784 561430 596840
rect 561498 596784 561554 596840
rect 561622 596784 561678 596840
rect 561250 580294 561306 580350
rect 561374 580294 561430 580350
rect 561498 580294 561554 580350
rect 561622 580294 561678 580350
rect 561250 580170 561306 580226
rect 561374 580170 561430 580226
rect 561498 580170 561554 580226
rect 561622 580170 561678 580226
rect 561250 580046 561306 580102
rect 561374 580046 561430 580102
rect 561498 580046 561554 580102
rect 561622 580046 561678 580102
rect 561250 579922 561306 579978
rect 561374 579922 561430 579978
rect 561498 579922 561554 579978
rect 561622 579922 561678 579978
rect 561250 562294 561306 562350
rect 561374 562294 561430 562350
rect 561498 562294 561554 562350
rect 561622 562294 561678 562350
rect 561250 562170 561306 562226
rect 561374 562170 561430 562226
rect 561498 562170 561554 562226
rect 561622 562170 561678 562226
rect 561250 562046 561306 562102
rect 561374 562046 561430 562102
rect 561498 562046 561554 562102
rect 561622 562046 561678 562102
rect 561250 561922 561306 561978
rect 561374 561922 561430 561978
rect 561498 561922 561554 561978
rect 561622 561922 561678 561978
rect 561250 544294 561306 544350
rect 561374 544294 561430 544350
rect 561498 544294 561554 544350
rect 561622 544294 561678 544350
rect 561250 544170 561306 544226
rect 561374 544170 561430 544226
rect 561498 544170 561554 544226
rect 561622 544170 561678 544226
rect 561250 544046 561306 544102
rect 561374 544046 561430 544102
rect 561498 544046 561554 544102
rect 561622 544046 561678 544102
rect 561250 543922 561306 543978
rect 561374 543922 561430 543978
rect 561498 543922 561554 543978
rect 561622 543922 561678 543978
rect 111250 526294 111306 526350
rect 111374 526294 111430 526350
rect 111498 526294 111554 526350
rect 111622 526294 111678 526350
rect 111250 526170 111306 526226
rect 111374 526170 111430 526226
rect 111498 526170 111554 526226
rect 111622 526170 111678 526226
rect 111250 526046 111306 526102
rect 111374 526046 111430 526102
rect 111498 526046 111554 526102
rect 111622 526046 111678 526102
rect 111250 525922 111306 525978
rect 111374 525922 111430 525978
rect 111498 525922 111554 525978
rect 111622 525922 111678 525978
rect 96970 514294 97026 514350
rect 97094 514294 97150 514350
rect 97218 514294 97274 514350
rect 97342 514294 97398 514350
rect 96970 514170 97026 514226
rect 97094 514170 97150 514226
rect 97218 514170 97274 514226
rect 97342 514170 97398 514226
rect 96970 514046 97026 514102
rect 97094 514046 97150 514102
rect 97218 514046 97274 514102
rect 97342 514046 97398 514102
rect 96970 513922 97026 513978
rect 97094 513922 97150 513978
rect 97218 513922 97274 513978
rect 97342 513922 97398 513978
rect 100598 514294 100654 514350
rect 100722 514294 100778 514350
rect 100598 514170 100654 514226
rect 100722 514170 100778 514226
rect 100598 514046 100654 514102
rect 100722 514046 100778 514102
rect 100598 513922 100654 513978
rect 100722 513922 100778 513978
rect 115958 526237 116014 526293
rect 116082 526237 116138 526293
rect 115958 526113 116014 526169
rect 116082 526113 116138 526169
rect 115958 525989 116014 526045
rect 116082 525989 116138 526045
rect 115958 525865 116014 525921
rect 116082 525865 116138 525921
rect 146678 526237 146734 526293
rect 146802 526237 146858 526293
rect 146678 526113 146734 526169
rect 146802 526113 146858 526169
rect 146678 525989 146734 526045
rect 146802 525989 146858 526045
rect 146678 525865 146734 525921
rect 146802 525865 146858 525921
rect 177398 526237 177454 526293
rect 177522 526237 177578 526293
rect 177398 526113 177454 526169
rect 177522 526113 177578 526169
rect 177398 525989 177454 526045
rect 177522 525989 177578 526045
rect 177398 525865 177454 525921
rect 177522 525865 177578 525921
rect 208118 526237 208174 526293
rect 208242 526237 208298 526293
rect 208118 526113 208174 526169
rect 208242 526113 208298 526169
rect 208118 525989 208174 526045
rect 208242 525989 208298 526045
rect 208118 525865 208174 525921
rect 208242 525865 208298 525921
rect 238838 526237 238894 526293
rect 238962 526237 239018 526293
rect 238838 526113 238894 526169
rect 238962 526113 239018 526169
rect 238838 525989 238894 526045
rect 238962 525989 239018 526045
rect 238838 525865 238894 525921
rect 238962 525865 239018 525921
rect 269558 526237 269614 526293
rect 269682 526237 269738 526293
rect 269558 526113 269614 526169
rect 269682 526113 269738 526169
rect 269558 525989 269614 526045
rect 269682 525989 269738 526045
rect 269558 525865 269614 525921
rect 269682 525865 269738 525921
rect 300278 526237 300334 526293
rect 300402 526237 300458 526293
rect 300278 526113 300334 526169
rect 300402 526113 300458 526169
rect 300278 525989 300334 526045
rect 300402 525989 300458 526045
rect 300278 525865 300334 525921
rect 300402 525865 300458 525921
rect 330998 526237 331054 526293
rect 331122 526237 331178 526293
rect 330998 526113 331054 526169
rect 331122 526113 331178 526169
rect 330998 525989 331054 526045
rect 331122 525989 331178 526045
rect 330998 525865 331054 525921
rect 331122 525865 331178 525921
rect 361718 526237 361774 526293
rect 361842 526237 361898 526293
rect 361718 526113 361774 526169
rect 361842 526113 361898 526169
rect 361718 525989 361774 526045
rect 361842 525989 361898 526045
rect 361718 525865 361774 525921
rect 361842 525865 361898 525921
rect 392438 526237 392494 526293
rect 392562 526237 392618 526293
rect 392438 526113 392494 526169
rect 392562 526113 392618 526169
rect 392438 525989 392494 526045
rect 392562 525989 392618 526045
rect 392438 525865 392494 525921
rect 392562 525865 392618 525921
rect 423158 526237 423214 526293
rect 423282 526237 423338 526293
rect 423158 526113 423214 526169
rect 423282 526113 423338 526169
rect 423158 525989 423214 526045
rect 423282 525989 423338 526045
rect 423158 525865 423214 525921
rect 423282 525865 423338 525921
rect 453878 526237 453934 526293
rect 454002 526237 454058 526293
rect 453878 526113 453934 526169
rect 454002 526113 454058 526169
rect 453878 525989 453934 526045
rect 454002 525989 454058 526045
rect 453878 525865 453934 525921
rect 454002 525865 454058 525921
rect 484598 526237 484654 526293
rect 484722 526237 484778 526293
rect 484598 526113 484654 526169
rect 484722 526113 484778 526169
rect 484598 525989 484654 526045
rect 484722 525989 484778 526045
rect 484598 525865 484654 525921
rect 484722 525865 484778 525921
rect 515318 526237 515374 526293
rect 515442 526237 515498 526293
rect 515318 526113 515374 526169
rect 515442 526113 515498 526169
rect 515318 525989 515374 526045
rect 515442 525989 515498 526045
rect 515318 525865 515374 525921
rect 515442 525865 515498 525921
rect 546038 526237 546094 526293
rect 546162 526237 546218 526293
rect 546038 526113 546094 526169
rect 546162 526113 546218 526169
rect 546038 525989 546094 526045
rect 546162 525989 546218 526045
rect 546038 525865 546094 525921
rect 546162 525865 546218 525921
rect 561250 526294 561306 526350
rect 561374 526294 561430 526350
rect 561498 526294 561554 526350
rect 561622 526294 561678 526350
rect 561250 526170 561306 526226
rect 561374 526170 561430 526226
rect 561498 526170 561554 526226
rect 561622 526170 561678 526226
rect 561250 526046 561306 526102
rect 561374 526046 561430 526102
rect 561498 526046 561554 526102
rect 561622 526046 561678 526102
rect 561250 525922 561306 525978
rect 561374 525922 561430 525978
rect 561498 525922 561554 525978
rect 561622 525922 561678 525978
rect 131318 514294 131374 514350
rect 131442 514294 131498 514350
rect 131318 514170 131374 514226
rect 131442 514170 131498 514226
rect 131318 514046 131374 514102
rect 131442 514046 131498 514102
rect 131318 513922 131374 513978
rect 131442 513922 131498 513978
rect 162038 514294 162094 514350
rect 162162 514294 162218 514350
rect 162038 514170 162094 514226
rect 162162 514170 162218 514226
rect 162038 514046 162094 514102
rect 162162 514046 162218 514102
rect 162038 513922 162094 513978
rect 162162 513922 162218 513978
rect 192758 514294 192814 514350
rect 192882 514294 192938 514350
rect 192758 514170 192814 514226
rect 192882 514170 192938 514226
rect 192758 514046 192814 514102
rect 192882 514046 192938 514102
rect 192758 513922 192814 513978
rect 192882 513922 192938 513978
rect 223478 514294 223534 514350
rect 223602 514294 223658 514350
rect 223478 514170 223534 514226
rect 223602 514170 223658 514226
rect 223478 514046 223534 514102
rect 223602 514046 223658 514102
rect 223478 513922 223534 513978
rect 223602 513922 223658 513978
rect 254198 514294 254254 514350
rect 254322 514294 254378 514350
rect 254198 514170 254254 514226
rect 254322 514170 254378 514226
rect 254198 514046 254254 514102
rect 254322 514046 254378 514102
rect 254198 513922 254254 513978
rect 254322 513922 254378 513978
rect 284918 514294 284974 514350
rect 285042 514294 285098 514350
rect 284918 514170 284974 514226
rect 285042 514170 285098 514226
rect 284918 514046 284974 514102
rect 285042 514046 285098 514102
rect 284918 513922 284974 513978
rect 285042 513922 285098 513978
rect 315638 514294 315694 514350
rect 315762 514294 315818 514350
rect 315638 514170 315694 514226
rect 315762 514170 315818 514226
rect 315638 514046 315694 514102
rect 315762 514046 315818 514102
rect 315638 513922 315694 513978
rect 315762 513922 315818 513978
rect 346358 514294 346414 514350
rect 346482 514294 346538 514350
rect 346358 514170 346414 514226
rect 346482 514170 346538 514226
rect 346358 514046 346414 514102
rect 346482 514046 346538 514102
rect 346358 513922 346414 513978
rect 346482 513922 346538 513978
rect 377078 514294 377134 514350
rect 377202 514294 377258 514350
rect 377078 514170 377134 514226
rect 377202 514170 377258 514226
rect 377078 514046 377134 514102
rect 377202 514046 377258 514102
rect 377078 513922 377134 513978
rect 377202 513922 377258 513978
rect 407798 514294 407854 514350
rect 407922 514294 407978 514350
rect 407798 514170 407854 514226
rect 407922 514170 407978 514226
rect 407798 514046 407854 514102
rect 407922 514046 407978 514102
rect 407798 513922 407854 513978
rect 407922 513922 407978 513978
rect 438518 514294 438574 514350
rect 438642 514294 438698 514350
rect 438518 514170 438574 514226
rect 438642 514170 438698 514226
rect 438518 514046 438574 514102
rect 438642 514046 438698 514102
rect 438518 513922 438574 513978
rect 438642 513922 438698 513978
rect 469238 514294 469294 514350
rect 469362 514294 469418 514350
rect 469238 514170 469294 514226
rect 469362 514170 469418 514226
rect 469238 514046 469294 514102
rect 469362 514046 469418 514102
rect 469238 513922 469294 513978
rect 469362 513922 469418 513978
rect 499958 514294 500014 514350
rect 500082 514294 500138 514350
rect 499958 514170 500014 514226
rect 500082 514170 500138 514226
rect 499958 514046 500014 514102
rect 500082 514046 500138 514102
rect 499958 513922 500014 513978
rect 500082 513922 500138 513978
rect 530678 514294 530734 514350
rect 530802 514294 530858 514350
rect 530678 514170 530734 514226
rect 530802 514170 530858 514226
rect 530678 514046 530734 514102
rect 530802 514046 530858 514102
rect 530678 513922 530734 513978
rect 530802 513922 530858 513978
rect 111250 508294 111306 508350
rect 111374 508294 111430 508350
rect 111498 508294 111554 508350
rect 111622 508294 111678 508350
rect 111250 508170 111306 508226
rect 111374 508170 111430 508226
rect 111498 508170 111554 508226
rect 111622 508170 111678 508226
rect 111250 508046 111306 508102
rect 111374 508046 111430 508102
rect 111498 508046 111554 508102
rect 111622 508046 111678 508102
rect 111250 507922 111306 507978
rect 111374 507922 111430 507978
rect 111498 507922 111554 507978
rect 111622 507922 111678 507978
rect 96970 496294 97026 496350
rect 97094 496294 97150 496350
rect 97218 496294 97274 496350
rect 97342 496294 97398 496350
rect 96970 496170 97026 496226
rect 97094 496170 97150 496226
rect 97218 496170 97274 496226
rect 97342 496170 97398 496226
rect 96970 496046 97026 496102
rect 97094 496046 97150 496102
rect 97218 496046 97274 496102
rect 97342 496046 97398 496102
rect 96970 495922 97026 495978
rect 97094 495922 97150 495978
rect 97218 495922 97274 495978
rect 97342 495922 97398 495978
rect 100598 496294 100654 496350
rect 100722 496294 100778 496350
rect 100598 496170 100654 496226
rect 100722 496170 100778 496226
rect 100598 496046 100654 496102
rect 100722 496046 100778 496102
rect 100598 495922 100654 495978
rect 100722 495922 100778 495978
rect 115958 508294 116014 508350
rect 116082 508294 116138 508350
rect 115958 508170 116014 508226
rect 116082 508170 116138 508226
rect 115958 508046 116014 508102
rect 116082 508046 116138 508102
rect 115958 507922 116014 507978
rect 116082 507922 116138 507978
rect 146678 508294 146734 508350
rect 146802 508294 146858 508350
rect 146678 508170 146734 508226
rect 146802 508170 146858 508226
rect 146678 508046 146734 508102
rect 146802 508046 146858 508102
rect 146678 507922 146734 507978
rect 146802 507922 146858 507978
rect 177398 508294 177454 508350
rect 177522 508294 177578 508350
rect 177398 508170 177454 508226
rect 177522 508170 177578 508226
rect 177398 508046 177454 508102
rect 177522 508046 177578 508102
rect 177398 507922 177454 507978
rect 177522 507922 177578 507978
rect 208118 508294 208174 508350
rect 208242 508294 208298 508350
rect 208118 508170 208174 508226
rect 208242 508170 208298 508226
rect 208118 508046 208174 508102
rect 208242 508046 208298 508102
rect 208118 507922 208174 507978
rect 208242 507922 208298 507978
rect 238838 508294 238894 508350
rect 238962 508294 239018 508350
rect 238838 508170 238894 508226
rect 238962 508170 239018 508226
rect 238838 508046 238894 508102
rect 238962 508046 239018 508102
rect 238838 507922 238894 507978
rect 238962 507922 239018 507978
rect 269558 508294 269614 508350
rect 269682 508294 269738 508350
rect 269558 508170 269614 508226
rect 269682 508170 269738 508226
rect 269558 508046 269614 508102
rect 269682 508046 269738 508102
rect 269558 507922 269614 507978
rect 269682 507922 269738 507978
rect 300278 508294 300334 508350
rect 300402 508294 300458 508350
rect 300278 508170 300334 508226
rect 300402 508170 300458 508226
rect 300278 508046 300334 508102
rect 300402 508046 300458 508102
rect 300278 507922 300334 507978
rect 300402 507922 300458 507978
rect 330998 508294 331054 508350
rect 331122 508294 331178 508350
rect 330998 508170 331054 508226
rect 331122 508170 331178 508226
rect 330998 508046 331054 508102
rect 331122 508046 331178 508102
rect 330998 507922 331054 507978
rect 331122 507922 331178 507978
rect 361718 508294 361774 508350
rect 361842 508294 361898 508350
rect 361718 508170 361774 508226
rect 361842 508170 361898 508226
rect 361718 508046 361774 508102
rect 361842 508046 361898 508102
rect 361718 507922 361774 507978
rect 361842 507922 361898 507978
rect 392438 508294 392494 508350
rect 392562 508294 392618 508350
rect 392438 508170 392494 508226
rect 392562 508170 392618 508226
rect 392438 508046 392494 508102
rect 392562 508046 392618 508102
rect 392438 507922 392494 507978
rect 392562 507922 392618 507978
rect 423158 508294 423214 508350
rect 423282 508294 423338 508350
rect 423158 508170 423214 508226
rect 423282 508170 423338 508226
rect 423158 508046 423214 508102
rect 423282 508046 423338 508102
rect 423158 507922 423214 507978
rect 423282 507922 423338 507978
rect 453878 508294 453934 508350
rect 454002 508294 454058 508350
rect 453878 508170 453934 508226
rect 454002 508170 454058 508226
rect 453878 508046 453934 508102
rect 454002 508046 454058 508102
rect 453878 507922 453934 507978
rect 454002 507922 454058 507978
rect 484598 508294 484654 508350
rect 484722 508294 484778 508350
rect 484598 508170 484654 508226
rect 484722 508170 484778 508226
rect 484598 508046 484654 508102
rect 484722 508046 484778 508102
rect 484598 507922 484654 507978
rect 484722 507922 484778 507978
rect 515318 508294 515374 508350
rect 515442 508294 515498 508350
rect 515318 508170 515374 508226
rect 515442 508170 515498 508226
rect 515318 508046 515374 508102
rect 515442 508046 515498 508102
rect 515318 507922 515374 507978
rect 515442 507922 515498 507978
rect 546038 508294 546094 508350
rect 546162 508294 546218 508350
rect 546038 508170 546094 508226
rect 546162 508170 546218 508226
rect 546038 508046 546094 508102
rect 546162 508046 546218 508102
rect 546038 507922 546094 507978
rect 546162 507922 546218 507978
rect 561250 508294 561306 508350
rect 561374 508294 561430 508350
rect 561498 508294 561554 508350
rect 561622 508294 561678 508350
rect 561250 508170 561306 508226
rect 561374 508170 561430 508226
rect 561498 508170 561554 508226
rect 561622 508170 561678 508226
rect 561250 508046 561306 508102
rect 561374 508046 561430 508102
rect 561498 508046 561554 508102
rect 561622 508046 561678 508102
rect 561250 507922 561306 507978
rect 561374 507922 561430 507978
rect 561498 507922 561554 507978
rect 561622 507922 561678 507978
rect 131318 496294 131374 496350
rect 131442 496294 131498 496350
rect 131318 496170 131374 496226
rect 131442 496170 131498 496226
rect 131318 496046 131374 496102
rect 131442 496046 131498 496102
rect 131318 495922 131374 495978
rect 131442 495922 131498 495978
rect 162038 496294 162094 496350
rect 162162 496294 162218 496350
rect 162038 496170 162094 496226
rect 162162 496170 162218 496226
rect 162038 496046 162094 496102
rect 162162 496046 162218 496102
rect 162038 495922 162094 495978
rect 162162 495922 162218 495978
rect 192758 496294 192814 496350
rect 192882 496294 192938 496350
rect 192758 496170 192814 496226
rect 192882 496170 192938 496226
rect 192758 496046 192814 496102
rect 192882 496046 192938 496102
rect 192758 495922 192814 495978
rect 192882 495922 192938 495978
rect 223478 496294 223534 496350
rect 223602 496294 223658 496350
rect 223478 496170 223534 496226
rect 223602 496170 223658 496226
rect 223478 496046 223534 496102
rect 223602 496046 223658 496102
rect 223478 495922 223534 495978
rect 223602 495922 223658 495978
rect 254198 496294 254254 496350
rect 254322 496294 254378 496350
rect 254198 496170 254254 496226
rect 254322 496170 254378 496226
rect 254198 496046 254254 496102
rect 254322 496046 254378 496102
rect 254198 495922 254254 495978
rect 254322 495922 254378 495978
rect 284918 496294 284974 496350
rect 285042 496294 285098 496350
rect 284918 496170 284974 496226
rect 285042 496170 285098 496226
rect 284918 496046 284974 496102
rect 285042 496046 285098 496102
rect 284918 495922 284974 495978
rect 285042 495922 285098 495978
rect 315638 496294 315694 496350
rect 315762 496294 315818 496350
rect 315638 496170 315694 496226
rect 315762 496170 315818 496226
rect 315638 496046 315694 496102
rect 315762 496046 315818 496102
rect 315638 495922 315694 495978
rect 315762 495922 315818 495978
rect 346358 496294 346414 496350
rect 346482 496294 346538 496350
rect 346358 496170 346414 496226
rect 346482 496170 346538 496226
rect 346358 496046 346414 496102
rect 346482 496046 346538 496102
rect 346358 495922 346414 495978
rect 346482 495922 346538 495978
rect 377078 496294 377134 496350
rect 377202 496294 377258 496350
rect 377078 496170 377134 496226
rect 377202 496170 377258 496226
rect 377078 496046 377134 496102
rect 377202 496046 377258 496102
rect 377078 495922 377134 495978
rect 377202 495922 377258 495978
rect 407798 496294 407854 496350
rect 407922 496294 407978 496350
rect 407798 496170 407854 496226
rect 407922 496170 407978 496226
rect 407798 496046 407854 496102
rect 407922 496046 407978 496102
rect 407798 495922 407854 495978
rect 407922 495922 407978 495978
rect 438518 496294 438574 496350
rect 438642 496294 438698 496350
rect 438518 496170 438574 496226
rect 438642 496170 438698 496226
rect 438518 496046 438574 496102
rect 438642 496046 438698 496102
rect 438518 495922 438574 495978
rect 438642 495922 438698 495978
rect 469238 496294 469294 496350
rect 469362 496294 469418 496350
rect 469238 496170 469294 496226
rect 469362 496170 469418 496226
rect 469238 496046 469294 496102
rect 469362 496046 469418 496102
rect 469238 495922 469294 495978
rect 469362 495922 469418 495978
rect 499958 496294 500014 496350
rect 500082 496294 500138 496350
rect 499958 496170 500014 496226
rect 500082 496170 500138 496226
rect 499958 496046 500014 496102
rect 500082 496046 500138 496102
rect 499958 495922 500014 495978
rect 500082 495922 500138 495978
rect 530678 496294 530734 496350
rect 530802 496294 530858 496350
rect 530678 496170 530734 496226
rect 530802 496170 530858 496226
rect 530678 496046 530734 496102
rect 530802 496046 530858 496102
rect 530678 495922 530734 495978
rect 530802 495922 530858 495978
rect 111250 490294 111306 490350
rect 111374 490294 111430 490350
rect 111498 490294 111554 490350
rect 111622 490294 111678 490350
rect 111250 490170 111306 490226
rect 111374 490170 111430 490226
rect 111498 490170 111554 490226
rect 111622 490170 111678 490226
rect 111250 490046 111306 490102
rect 111374 490046 111430 490102
rect 111498 490046 111554 490102
rect 111622 490046 111678 490102
rect 111250 489922 111306 489978
rect 111374 489922 111430 489978
rect 111498 489922 111554 489978
rect 111622 489922 111678 489978
rect 96970 478294 97026 478350
rect 97094 478294 97150 478350
rect 97218 478294 97274 478350
rect 97342 478294 97398 478350
rect 96970 478170 97026 478226
rect 97094 478170 97150 478226
rect 97218 478170 97274 478226
rect 97342 478170 97398 478226
rect 96970 478046 97026 478102
rect 97094 478046 97150 478102
rect 97218 478046 97274 478102
rect 97342 478046 97398 478102
rect 96970 477922 97026 477978
rect 97094 477922 97150 477978
rect 97218 477922 97274 477978
rect 97342 477922 97398 477978
rect 100598 478294 100654 478350
rect 100722 478294 100778 478350
rect 100598 478170 100654 478226
rect 100722 478170 100778 478226
rect 100598 478046 100654 478102
rect 100722 478046 100778 478102
rect 100598 477922 100654 477978
rect 100722 477922 100778 477978
rect 115958 490294 116014 490350
rect 116082 490294 116138 490350
rect 115958 490170 116014 490226
rect 116082 490170 116138 490226
rect 115958 490046 116014 490102
rect 116082 490046 116138 490102
rect 115958 489922 116014 489978
rect 116082 489922 116138 489978
rect 146678 490294 146734 490350
rect 146802 490294 146858 490350
rect 146678 490170 146734 490226
rect 146802 490170 146858 490226
rect 146678 490046 146734 490102
rect 146802 490046 146858 490102
rect 146678 489922 146734 489978
rect 146802 489922 146858 489978
rect 177398 490294 177454 490350
rect 177522 490294 177578 490350
rect 177398 490170 177454 490226
rect 177522 490170 177578 490226
rect 177398 490046 177454 490102
rect 177522 490046 177578 490102
rect 177398 489922 177454 489978
rect 177522 489922 177578 489978
rect 208118 490294 208174 490350
rect 208242 490294 208298 490350
rect 208118 490170 208174 490226
rect 208242 490170 208298 490226
rect 208118 490046 208174 490102
rect 208242 490046 208298 490102
rect 208118 489922 208174 489978
rect 208242 489922 208298 489978
rect 238838 490294 238894 490350
rect 238962 490294 239018 490350
rect 238838 490170 238894 490226
rect 238962 490170 239018 490226
rect 238838 490046 238894 490102
rect 238962 490046 239018 490102
rect 238838 489922 238894 489978
rect 238962 489922 239018 489978
rect 269558 490294 269614 490350
rect 269682 490294 269738 490350
rect 269558 490170 269614 490226
rect 269682 490170 269738 490226
rect 269558 490046 269614 490102
rect 269682 490046 269738 490102
rect 269558 489922 269614 489978
rect 269682 489922 269738 489978
rect 300278 490294 300334 490350
rect 300402 490294 300458 490350
rect 300278 490170 300334 490226
rect 300402 490170 300458 490226
rect 300278 490046 300334 490102
rect 300402 490046 300458 490102
rect 300278 489922 300334 489978
rect 300402 489922 300458 489978
rect 330998 490294 331054 490350
rect 331122 490294 331178 490350
rect 330998 490170 331054 490226
rect 331122 490170 331178 490226
rect 330998 490046 331054 490102
rect 331122 490046 331178 490102
rect 330998 489922 331054 489978
rect 331122 489922 331178 489978
rect 361718 490294 361774 490350
rect 361842 490294 361898 490350
rect 361718 490170 361774 490226
rect 361842 490170 361898 490226
rect 361718 490046 361774 490102
rect 361842 490046 361898 490102
rect 361718 489922 361774 489978
rect 361842 489922 361898 489978
rect 392438 490294 392494 490350
rect 392562 490294 392618 490350
rect 392438 490170 392494 490226
rect 392562 490170 392618 490226
rect 392438 490046 392494 490102
rect 392562 490046 392618 490102
rect 392438 489922 392494 489978
rect 392562 489922 392618 489978
rect 423158 490294 423214 490350
rect 423282 490294 423338 490350
rect 423158 490170 423214 490226
rect 423282 490170 423338 490226
rect 423158 490046 423214 490102
rect 423282 490046 423338 490102
rect 423158 489922 423214 489978
rect 423282 489922 423338 489978
rect 453878 490294 453934 490350
rect 454002 490294 454058 490350
rect 453878 490170 453934 490226
rect 454002 490170 454058 490226
rect 453878 490046 453934 490102
rect 454002 490046 454058 490102
rect 453878 489922 453934 489978
rect 454002 489922 454058 489978
rect 484598 490294 484654 490350
rect 484722 490294 484778 490350
rect 484598 490170 484654 490226
rect 484722 490170 484778 490226
rect 484598 490046 484654 490102
rect 484722 490046 484778 490102
rect 484598 489922 484654 489978
rect 484722 489922 484778 489978
rect 515318 490294 515374 490350
rect 515442 490294 515498 490350
rect 515318 490170 515374 490226
rect 515442 490170 515498 490226
rect 515318 490046 515374 490102
rect 515442 490046 515498 490102
rect 515318 489922 515374 489978
rect 515442 489922 515498 489978
rect 546038 490294 546094 490350
rect 546162 490294 546218 490350
rect 546038 490170 546094 490226
rect 546162 490170 546218 490226
rect 546038 490046 546094 490102
rect 546162 490046 546218 490102
rect 546038 489922 546094 489978
rect 546162 489922 546218 489978
rect 561250 490294 561306 490350
rect 561374 490294 561430 490350
rect 561498 490294 561554 490350
rect 561622 490294 561678 490350
rect 561250 490170 561306 490226
rect 561374 490170 561430 490226
rect 561498 490170 561554 490226
rect 561622 490170 561678 490226
rect 561250 490046 561306 490102
rect 561374 490046 561430 490102
rect 561498 490046 561554 490102
rect 561622 490046 561678 490102
rect 561250 489922 561306 489978
rect 561374 489922 561430 489978
rect 561498 489922 561554 489978
rect 561622 489922 561678 489978
rect 131318 478294 131374 478350
rect 131442 478294 131498 478350
rect 131318 478170 131374 478226
rect 131442 478170 131498 478226
rect 131318 478046 131374 478102
rect 131442 478046 131498 478102
rect 131318 477922 131374 477978
rect 131442 477922 131498 477978
rect 162038 478294 162094 478350
rect 162162 478294 162218 478350
rect 162038 478170 162094 478226
rect 162162 478170 162218 478226
rect 162038 478046 162094 478102
rect 162162 478046 162218 478102
rect 162038 477922 162094 477978
rect 162162 477922 162218 477978
rect 192758 478294 192814 478350
rect 192882 478294 192938 478350
rect 192758 478170 192814 478226
rect 192882 478170 192938 478226
rect 192758 478046 192814 478102
rect 192882 478046 192938 478102
rect 192758 477922 192814 477978
rect 192882 477922 192938 477978
rect 223478 478294 223534 478350
rect 223602 478294 223658 478350
rect 223478 478170 223534 478226
rect 223602 478170 223658 478226
rect 223478 478046 223534 478102
rect 223602 478046 223658 478102
rect 223478 477922 223534 477978
rect 223602 477922 223658 477978
rect 254198 478294 254254 478350
rect 254322 478294 254378 478350
rect 254198 478170 254254 478226
rect 254322 478170 254378 478226
rect 254198 478046 254254 478102
rect 254322 478046 254378 478102
rect 254198 477922 254254 477978
rect 254322 477922 254378 477978
rect 284918 478294 284974 478350
rect 285042 478294 285098 478350
rect 284918 478170 284974 478226
rect 285042 478170 285098 478226
rect 284918 478046 284974 478102
rect 285042 478046 285098 478102
rect 284918 477922 284974 477978
rect 285042 477922 285098 477978
rect 315638 478294 315694 478350
rect 315762 478294 315818 478350
rect 315638 478170 315694 478226
rect 315762 478170 315818 478226
rect 315638 478046 315694 478102
rect 315762 478046 315818 478102
rect 315638 477922 315694 477978
rect 315762 477922 315818 477978
rect 346358 478294 346414 478350
rect 346482 478294 346538 478350
rect 346358 478170 346414 478226
rect 346482 478170 346538 478226
rect 346358 478046 346414 478102
rect 346482 478046 346538 478102
rect 346358 477922 346414 477978
rect 346482 477922 346538 477978
rect 377078 478294 377134 478350
rect 377202 478294 377258 478350
rect 377078 478170 377134 478226
rect 377202 478170 377258 478226
rect 377078 478046 377134 478102
rect 377202 478046 377258 478102
rect 377078 477922 377134 477978
rect 377202 477922 377258 477978
rect 407798 478294 407854 478350
rect 407922 478294 407978 478350
rect 407798 478170 407854 478226
rect 407922 478170 407978 478226
rect 407798 478046 407854 478102
rect 407922 478046 407978 478102
rect 407798 477922 407854 477978
rect 407922 477922 407978 477978
rect 438518 478294 438574 478350
rect 438642 478294 438698 478350
rect 438518 478170 438574 478226
rect 438642 478170 438698 478226
rect 438518 478046 438574 478102
rect 438642 478046 438698 478102
rect 438518 477922 438574 477978
rect 438642 477922 438698 477978
rect 469238 478294 469294 478350
rect 469362 478294 469418 478350
rect 469238 478170 469294 478226
rect 469362 478170 469418 478226
rect 469238 478046 469294 478102
rect 469362 478046 469418 478102
rect 469238 477922 469294 477978
rect 469362 477922 469418 477978
rect 499958 478294 500014 478350
rect 500082 478294 500138 478350
rect 499958 478170 500014 478226
rect 500082 478170 500138 478226
rect 499958 478046 500014 478102
rect 500082 478046 500138 478102
rect 499958 477922 500014 477978
rect 500082 477922 500138 477978
rect 530678 478294 530734 478350
rect 530802 478294 530858 478350
rect 530678 478170 530734 478226
rect 530802 478170 530858 478226
rect 530678 478046 530734 478102
rect 530802 478046 530858 478102
rect 530678 477922 530734 477978
rect 530802 477922 530858 477978
rect 111250 472294 111306 472350
rect 111374 472294 111430 472350
rect 111498 472294 111554 472350
rect 111622 472294 111678 472350
rect 111250 472170 111306 472226
rect 111374 472170 111430 472226
rect 111498 472170 111554 472226
rect 111622 472170 111678 472226
rect 111250 472046 111306 472102
rect 111374 472046 111430 472102
rect 111498 472046 111554 472102
rect 111622 472046 111678 472102
rect 111250 471922 111306 471978
rect 111374 471922 111430 471978
rect 111498 471922 111554 471978
rect 111622 471922 111678 471978
rect 96970 460294 97026 460350
rect 97094 460294 97150 460350
rect 97218 460294 97274 460350
rect 97342 460294 97398 460350
rect 96970 460170 97026 460226
rect 97094 460170 97150 460226
rect 97218 460170 97274 460226
rect 97342 460170 97398 460226
rect 96970 460046 97026 460102
rect 97094 460046 97150 460102
rect 97218 460046 97274 460102
rect 97342 460046 97398 460102
rect 96970 459922 97026 459978
rect 97094 459922 97150 459978
rect 97218 459922 97274 459978
rect 97342 459922 97398 459978
rect 100598 460294 100654 460350
rect 100722 460294 100778 460350
rect 100598 460170 100654 460226
rect 100722 460170 100778 460226
rect 100598 460046 100654 460102
rect 100722 460046 100778 460102
rect 100598 459922 100654 459978
rect 100722 459922 100778 459978
rect 115958 472294 116014 472350
rect 116082 472294 116138 472350
rect 115958 472170 116014 472226
rect 116082 472170 116138 472226
rect 115958 472046 116014 472102
rect 116082 472046 116138 472102
rect 115958 471922 116014 471978
rect 116082 471922 116138 471978
rect 146678 472294 146734 472350
rect 146802 472294 146858 472350
rect 146678 472170 146734 472226
rect 146802 472170 146858 472226
rect 146678 472046 146734 472102
rect 146802 472046 146858 472102
rect 146678 471922 146734 471978
rect 146802 471922 146858 471978
rect 177398 472294 177454 472350
rect 177522 472294 177578 472350
rect 177398 472170 177454 472226
rect 177522 472170 177578 472226
rect 177398 472046 177454 472102
rect 177522 472046 177578 472102
rect 177398 471922 177454 471978
rect 177522 471922 177578 471978
rect 208118 472294 208174 472350
rect 208242 472294 208298 472350
rect 208118 472170 208174 472226
rect 208242 472170 208298 472226
rect 208118 472046 208174 472102
rect 208242 472046 208298 472102
rect 208118 471922 208174 471978
rect 208242 471922 208298 471978
rect 238838 472294 238894 472350
rect 238962 472294 239018 472350
rect 238838 472170 238894 472226
rect 238962 472170 239018 472226
rect 238838 472046 238894 472102
rect 238962 472046 239018 472102
rect 238838 471922 238894 471978
rect 238962 471922 239018 471978
rect 269558 472294 269614 472350
rect 269682 472294 269738 472350
rect 269558 472170 269614 472226
rect 269682 472170 269738 472226
rect 269558 472046 269614 472102
rect 269682 472046 269738 472102
rect 269558 471922 269614 471978
rect 269682 471922 269738 471978
rect 300278 472294 300334 472350
rect 300402 472294 300458 472350
rect 300278 472170 300334 472226
rect 300402 472170 300458 472226
rect 300278 472046 300334 472102
rect 300402 472046 300458 472102
rect 300278 471922 300334 471978
rect 300402 471922 300458 471978
rect 330998 472294 331054 472350
rect 331122 472294 331178 472350
rect 330998 472170 331054 472226
rect 331122 472170 331178 472226
rect 330998 472046 331054 472102
rect 331122 472046 331178 472102
rect 330998 471922 331054 471978
rect 331122 471922 331178 471978
rect 361718 472294 361774 472350
rect 361842 472294 361898 472350
rect 361718 472170 361774 472226
rect 361842 472170 361898 472226
rect 361718 472046 361774 472102
rect 361842 472046 361898 472102
rect 361718 471922 361774 471978
rect 361842 471922 361898 471978
rect 392438 472294 392494 472350
rect 392562 472294 392618 472350
rect 392438 472170 392494 472226
rect 392562 472170 392618 472226
rect 392438 472046 392494 472102
rect 392562 472046 392618 472102
rect 392438 471922 392494 471978
rect 392562 471922 392618 471978
rect 423158 472294 423214 472350
rect 423282 472294 423338 472350
rect 423158 472170 423214 472226
rect 423282 472170 423338 472226
rect 423158 472046 423214 472102
rect 423282 472046 423338 472102
rect 423158 471922 423214 471978
rect 423282 471922 423338 471978
rect 453878 472294 453934 472350
rect 454002 472294 454058 472350
rect 453878 472170 453934 472226
rect 454002 472170 454058 472226
rect 453878 472046 453934 472102
rect 454002 472046 454058 472102
rect 453878 471922 453934 471978
rect 454002 471922 454058 471978
rect 484598 472294 484654 472350
rect 484722 472294 484778 472350
rect 484598 472170 484654 472226
rect 484722 472170 484778 472226
rect 484598 472046 484654 472102
rect 484722 472046 484778 472102
rect 484598 471922 484654 471978
rect 484722 471922 484778 471978
rect 515318 472294 515374 472350
rect 515442 472294 515498 472350
rect 515318 472170 515374 472226
rect 515442 472170 515498 472226
rect 515318 472046 515374 472102
rect 515442 472046 515498 472102
rect 515318 471922 515374 471978
rect 515442 471922 515498 471978
rect 546038 472294 546094 472350
rect 546162 472294 546218 472350
rect 546038 472170 546094 472226
rect 546162 472170 546218 472226
rect 546038 472046 546094 472102
rect 546162 472046 546218 472102
rect 546038 471922 546094 471978
rect 546162 471922 546218 471978
rect 561250 472294 561306 472350
rect 561374 472294 561430 472350
rect 561498 472294 561554 472350
rect 561622 472294 561678 472350
rect 561250 472170 561306 472226
rect 561374 472170 561430 472226
rect 561498 472170 561554 472226
rect 561622 472170 561678 472226
rect 561250 472046 561306 472102
rect 561374 472046 561430 472102
rect 561498 472046 561554 472102
rect 561622 472046 561678 472102
rect 561250 471922 561306 471978
rect 561374 471922 561430 471978
rect 561498 471922 561554 471978
rect 561622 471922 561678 471978
rect 131318 460294 131374 460350
rect 131442 460294 131498 460350
rect 131318 460170 131374 460226
rect 131442 460170 131498 460226
rect 131318 460046 131374 460102
rect 131442 460046 131498 460102
rect 131318 459922 131374 459978
rect 131442 459922 131498 459978
rect 162038 460294 162094 460350
rect 162162 460294 162218 460350
rect 162038 460170 162094 460226
rect 162162 460170 162218 460226
rect 162038 460046 162094 460102
rect 162162 460046 162218 460102
rect 162038 459922 162094 459978
rect 162162 459922 162218 459978
rect 192758 460294 192814 460350
rect 192882 460294 192938 460350
rect 192758 460170 192814 460226
rect 192882 460170 192938 460226
rect 192758 460046 192814 460102
rect 192882 460046 192938 460102
rect 192758 459922 192814 459978
rect 192882 459922 192938 459978
rect 223478 460294 223534 460350
rect 223602 460294 223658 460350
rect 223478 460170 223534 460226
rect 223602 460170 223658 460226
rect 223478 460046 223534 460102
rect 223602 460046 223658 460102
rect 223478 459922 223534 459978
rect 223602 459922 223658 459978
rect 254198 460294 254254 460350
rect 254322 460294 254378 460350
rect 254198 460170 254254 460226
rect 254322 460170 254378 460226
rect 254198 460046 254254 460102
rect 254322 460046 254378 460102
rect 254198 459922 254254 459978
rect 254322 459922 254378 459978
rect 284918 460294 284974 460350
rect 285042 460294 285098 460350
rect 284918 460170 284974 460226
rect 285042 460170 285098 460226
rect 284918 460046 284974 460102
rect 285042 460046 285098 460102
rect 284918 459922 284974 459978
rect 285042 459922 285098 459978
rect 315638 460294 315694 460350
rect 315762 460294 315818 460350
rect 315638 460170 315694 460226
rect 315762 460170 315818 460226
rect 315638 460046 315694 460102
rect 315762 460046 315818 460102
rect 315638 459922 315694 459978
rect 315762 459922 315818 459978
rect 346358 460294 346414 460350
rect 346482 460294 346538 460350
rect 346358 460170 346414 460226
rect 346482 460170 346538 460226
rect 346358 460046 346414 460102
rect 346482 460046 346538 460102
rect 346358 459922 346414 459978
rect 346482 459922 346538 459978
rect 377078 460294 377134 460350
rect 377202 460294 377258 460350
rect 377078 460170 377134 460226
rect 377202 460170 377258 460226
rect 377078 460046 377134 460102
rect 377202 460046 377258 460102
rect 377078 459922 377134 459978
rect 377202 459922 377258 459978
rect 407798 460294 407854 460350
rect 407922 460294 407978 460350
rect 407798 460170 407854 460226
rect 407922 460170 407978 460226
rect 407798 460046 407854 460102
rect 407922 460046 407978 460102
rect 407798 459922 407854 459978
rect 407922 459922 407978 459978
rect 438518 460294 438574 460350
rect 438642 460294 438698 460350
rect 438518 460170 438574 460226
rect 438642 460170 438698 460226
rect 438518 460046 438574 460102
rect 438642 460046 438698 460102
rect 438518 459922 438574 459978
rect 438642 459922 438698 459978
rect 469238 460294 469294 460350
rect 469362 460294 469418 460350
rect 469238 460170 469294 460226
rect 469362 460170 469418 460226
rect 469238 460046 469294 460102
rect 469362 460046 469418 460102
rect 469238 459922 469294 459978
rect 469362 459922 469418 459978
rect 499958 460294 500014 460350
rect 500082 460294 500138 460350
rect 499958 460170 500014 460226
rect 500082 460170 500138 460226
rect 499958 460046 500014 460102
rect 500082 460046 500138 460102
rect 499958 459922 500014 459978
rect 500082 459922 500138 459978
rect 530678 460294 530734 460350
rect 530802 460294 530858 460350
rect 530678 460170 530734 460226
rect 530802 460170 530858 460226
rect 530678 460046 530734 460102
rect 530802 460046 530858 460102
rect 530678 459922 530734 459978
rect 530802 459922 530858 459978
rect 111250 454294 111306 454350
rect 111374 454294 111430 454350
rect 111498 454294 111554 454350
rect 111622 454294 111678 454350
rect 111250 454170 111306 454226
rect 111374 454170 111430 454226
rect 111498 454170 111554 454226
rect 111622 454170 111678 454226
rect 111250 454046 111306 454102
rect 111374 454046 111430 454102
rect 111498 454046 111554 454102
rect 111622 454046 111678 454102
rect 111250 453922 111306 453978
rect 111374 453922 111430 453978
rect 111498 453922 111554 453978
rect 111622 453922 111678 453978
rect 96970 442294 97026 442350
rect 97094 442294 97150 442350
rect 97218 442294 97274 442350
rect 97342 442294 97398 442350
rect 96970 442170 97026 442226
rect 97094 442170 97150 442226
rect 97218 442170 97274 442226
rect 97342 442170 97398 442226
rect 96970 442046 97026 442102
rect 97094 442046 97150 442102
rect 97218 442046 97274 442102
rect 97342 442046 97398 442102
rect 96970 441922 97026 441978
rect 97094 441922 97150 441978
rect 97218 441922 97274 441978
rect 97342 441922 97398 441978
rect 100598 442294 100654 442350
rect 100722 442294 100778 442350
rect 100598 442170 100654 442226
rect 100722 442170 100778 442226
rect 100598 442046 100654 442102
rect 100722 442046 100778 442102
rect 100598 441922 100654 441978
rect 100722 441922 100778 441978
rect 115958 454294 116014 454350
rect 116082 454294 116138 454350
rect 115958 454170 116014 454226
rect 116082 454170 116138 454226
rect 115958 454046 116014 454102
rect 116082 454046 116138 454102
rect 115958 453922 116014 453978
rect 116082 453922 116138 453978
rect 146678 454294 146734 454350
rect 146802 454294 146858 454350
rect 146678 454170 146734 454226
rect 146802 454170 146858 454226
rect 146678 454046 146734 454102
rect 146802 454046 146858 454102
rect 146678 453922 146734 453978
rect 146802 453922 146858 453978
rect 177398 454294 177454 454350
rect 177522 454294 177578 454350
rect 177398 454170 177454 454226
rect 177522 454170 177578 454226
rect 177398 454046 177454 454102
rect 177522 454046 177578 454102
rect 177398 453922 177454 453978
rect 177522 453922 177578 453978
rect 208118 454294 208174 454350
rect 208242 454294 208298 454350
rect 208118 454170 208174 454226
rect 208242 454170 208298 454226
rect 208118 454046 208174 454102
rect 208242 454046 208298 454102
rect 208118 453922 208174 453978
rect 208242 453922 208298 453978
rect 238838 454294 238894 454350
rect 238962 454294 239018 454350
rect 238838 454170 238894 454226
rect 238962 454170 239018 454226
rect 238838 454046 238894 454102
rect 238962 454046 239018 454102
rect 238838 453922 238894 453978
rect 238962 453922 239018 453978
rect 269558 454294 269614 454350
rect 269682 454294 269738 454350
rect 269558 454170 269614 454226
rect 269682 454170 269738 454226
rect 269558 454046 269614 454102
rect 269682 454046 269738 454102
rect 269558 453922 269614 453978
rect 269682 453922 269738 453978
rect 300278 454294 300334 454350
rect 300402 454294 300458 454350
rect 300278 454170 300334 454226
rect 300402 454170 300458 454226
rect 300278 454046 300334 454102
rect 300402 454046 300458 454102
rect 300278 453922 300334 453978
rect 300402 453922 300458 453978
rect 330998 454294 331054 454350
rect 331122 454294 331178 454350
rect 330998 454170 331054 454226
rect 331122 454170 331178 454226
rect 330998 454046 331054 454102
rect 331122 454046 331178 454102
rect 330998 453922 331054 453978
rect 331122 453922 331178 453978
rect 361718 454294 361774 454350
rect 361842 454294 361898 454350
rect 361718 454170 361774 454226
rect 361842 454170 361898 454226
rect 361718 454046 361774 454102
rect 361842 454046 361898 454102
rect 361718 453922 361774 453978
rect 361842 453922 361898 453978
rect 392438 454294 392494 454350
rect 392562 454294 392618 454350
rect 392438 454170 392494 454226
rect 392562 454170 392618 454226
rect 392438 454046 392494 454102
rect 392562 454046 392618 454102
rect 392438 453922 392494 453978
rect 392562 453922 392618 453978
rect 423158 454294 423214 454350
rect 423282 454294 423338 454350
rect 423158 454170 423214 454226
rect 423282 454170 423338 454226
rect 423158 454046 423214 454102
rect 423282 454046 423338 454102
rect 423158 453922 423214 453978
rect 423282 453922 423338 453978
rect 453878 454294 453934 454350
rect 454002 454294 454058 454350
rect 453878 454170 453934 454226
rect 454002 454170 454058 454226
rect 453878 454046 453934 454102
rect 454002 454046 454058 454102
rect 453878 453922 453934 453978
rect 454002 453922 454058 453978
rect 484598 454294 484654 454350
rect 484722 454294 484778 454350
rect 484598 454170 484654 454226
rect 484722 454170 484778 454226
rect 484598 454046 484654 454102
rect 484722 454046 484778 454102
rect 484598 453922 484654 453978
rect 484722 453922 484778 453978
rect 515318 454294 515374 454350
rect 515442 454294 515498 454350
rect 515318 454170 515374 454226
rect 515442 454170 515498 454226
rect 515318 454046 515374 454102
rect 515442 454046 515498 454102
rect 515318 453922 515374 453978
rect 515442 453922 515498 453978
rect 546038 454294 546094 454350
rect 546162 454294 546218 454350
rect 546038 454170 546094 454226
rect 546162 454170 546218 454226
rect 546038 454046 546094 454102
rect 546162 454046 546218 454102
rect 546038 453922 546094 453978
rect 546162 453922 546218 453978
rect 561250 454294 561306 454350
rect 561374 454294 561430 454350
rect 561498 454294 561554 454350
rect 561622 454294 561678 454350
rect 561250 454170 561306 454226
rect 561374 454170 561430 454226
rect 561498 454170 561554 454226
rect 561622 454170 561678 454226
rect 561250 454046 561306 454102
rect 561374 454046 561430 454102
rect 561498 454046 561554 454102
rect 561622 454046 561678 454102
rect 561250 453922 561306 453978
rect 561374 453922 561430 453978
rect 561498 453922 561554 453978
rect 561622 453922 561678 453978
rect 131318 442294 131374 442350
rect 131442 442294 131498 442350
rect 131318 442170 131374 442226
rect 131442 442170 131498 442226
rect 131318 442046 131374 442102
rect 131442 442046 131498 442102
rect 131318 441922 131374 441978
rect 131442 441922 131498 441978
rect 162038 442294 162094 442350
rect 162162 442294 162218 442350
rect 162038 442170 162094 442226
rect 162162 442170 162218 442226
rect 162038 442046 162094 442102
rect 162162 442046 162218 442102
rect 162038 441922 162094 441978
rect 162162 441922 162218 441978
rect 192758 442294 192814 442350
rect 192882 442294 192938 442350
rect 192758 442170 192814 442226
rect 192882 442170 192938 442226
rect 192758 442046 192814 442102
rect 192882 442046 192938 442102
rect 192758 441922 192814 441978
rect 192882 441922 192938 441978
rect 223478 442294 223534 442350
rect 223602 442294 223658 442350
rect 223478 442170 223534 442226
rect 223602 442170 223658 442226
rect 223478 442046 223534 442102
rect 223602 442046 223658 442102
rect 223478 441922 223534 441978
rect 223602 441922 223658 441978
rect 254198 442294 254254 442350
rect 254322 442294 254378 442350
rect 254198 442170 254254 442226
rect 254322 442170 254378 442226
rect 254198 442046 254254 442102
rect 254322 442046 254378 442102
rect 254198 441922 254254 441978
rect 254322 441922 254378 441978
rect 284918 442294 284974 442350
rect 285042 442294 285098 442350
rect 284918 442170 284974 442226
rect 285042 442170 285098 442226
rect 284918 442046 284974 442102
rect 285042 442046 285098 442102
rect 284918 441922 284974 441978
rect 285042 441922 285098 441978
rect 315638 442294 315694 442350
rect 315762 442294 315818 442350
rect 315638 442170 315694 442226
rect 315762 442170 315818 442226
rect 315638 442046 315694 442102
rect 315762 442046 315818 442102
rect 315638 441922 315694 441978
rect 315762 441922 315818 441978
rect 346358 442294 346414 442350
rect 346482 442294 346538 442350
rect 346358 442170 346414 442226
rect 346482 442170 346538 442226
rect 346358 442046 346414 442102
rect 346482 442046 346538 442102
rect 346358 441922 346414 441978
rect 346482 441922 346538 441978
rect 377078 442294 377134 442350
rect 377202 442294 377258 442350
rect 377078 442170 377134 442226
rect 377202 442170 377258 442226
rect 377078 442046 377134 442102
rect 377202 442046 377258 442102
rect 377078 441922 377134 441978
rect 377202 441922 377258 441978
rect 407798 442294 407854 442350
rect 407922 442294 407978 442350
rect 407798 442170 407854 442226
rect 407922 442170 407978 442226
rect 407798 442046 407854 442102
rect 407922 442046 407978 442102
rect 407798 441922 407854 441978
rect 407922 441922 407978 441978
rect 438518 442294 438574 442350
rect 438642 442294 438698 442350
rect 438518 442170 438574 442226
rect 438642 442170 438698 442226
rect 438518 442046 438574 442102
rect 438642 442046 438698 442102
rect 438518 441922 438574 441978
rect 438642 441922 438698 441978
rect 469238 442294 469294 442350
rect 469362 442294 469418 442350
rect 469238 442170 469294 442226
rect 469362 442170 469418 442226
rect 469238 442046 469294 442102
rect 469362 442046 469418 442102
rect 469238 441922 469294 441978
rect 469362 441922 469418 441978
rect 499958 442294 500014 442350
rect 500082 442294 500138 442350
rect 499958 442170 500014 442226
rect 500082 442170 500138 442226
rect 499958 442046 500014 442102
rect 500082 442046 500138 442102
rect 499958 441922 500014 441978
rect 500082 441922 500138 441978
rect 530678 442294 530734 442350
rect 530802 442294 530858 442350
rect 530678 442170 530734 442226
rect 530802 442170 530858 442226
rect 530678 442046 530734 442102
rect 530802 442046 530858 442102
rect 530678 441922 530734 441978
rect 530802 441922 530858 441978
rect 111250 436294 111306 436350
rect 111374 436294 111430 436350
rect 111498 436294 111554 436350
rect 111622 436294 111678 436350
rect 111250 436170 111306 436226
rect 111374 436170 111430 436226
rect 111498 436170 111554 436226
rect 111622 436170 111678 436226
rect 111250 436046 111306 436102
rect 111374 436046 111430 436102
rect 111498 436046 111554 436102
rect 111622 436046 111678 436102
rect 111250 435922 111306 435978
rect 111374 435922 111430 435978
rect 111498 435922 111554 435978
rect 111622 435922 111678 435978
rect 96970 424294 97026 424350
rect 97094 424294 97150 424350
rect 97218 424294 97274 424350
rect 97342 424294 97398 424350
rect 96970 424170 97026 424226
rect 97094 424170 97150 424226
rect 97218 424170 97274 424226
rect 97342 424170 97398 424226
rect 96970 424046 97026 424102
rect 97094 424046 97150 424102
rect 97218 424046 97274 424102
rect 97342 424046 97398 424102
rect 96970 423922 97026 423978
rect 97094 423922 97150 423978
rect 97218 423922 97274 423978
rect 97342 423922 97398 423978
rect 100598 424294 100654 424350
rect 100722 424294 100778 424350
rect 100598 424170 100654 424226
rect 100722 424170 100778 424226
rect 100598 424046 100654 424102
rect 100722 424046 100778 424102
rect 100598 423922 100654 423978
rect 100722 423922 100778 423978
rect 115958 436294 116014 436350
rect 116082 436294 116138 436350
rect 115958 436170 116014 436226
rect 116082 436170 116138 436226
rect 115958 436046 116014 436102
rect 116082 436046 116138 436102
rect 115958 435922 116014 435978
rect 116082 435922 116138 435978
rect 146678 436294 146734 436350
rect 146802 436294 146858 436350
rect 146678 436170 146734 436226
rect 146802 436170 146858 436226
rect 146678 436046 146734 436102
rect 146802 436046 146858 436102
rect 146678 435922 146734 435978
rect 146802 435922 146858 435978
rect 177398 436294 177454 436350
rect 177522 436294 177578 436350
rect 177398 436170 177454 436226
rect 177522 436170 177578 436226
rect 177398 436046 177454 436102
rect 177522 436046 177578 436102
rect 177398 435922 177454 435978
rect 177522 435922 177578 435978
rect 208118 436294 208174 436350
rect 208242 436294 208298 436350
rect 208118 436170 208174 436226
rect 208242 436170 208298 436226
rect 208118 436046 208174 436102
rect 208242 436046 208298 436102
rect 208118 435922 208174 435978
rect 208242 435922 208298 435978
rect 238838 436294 238894 436350
rect 238962 436294 239018 436350
rect 238838 436170 238894 436226
rect 238962 436170 239018 436226
rect 238838 436046 238894 436102
rect 238962 436046 239018 436102
rect 238838 435922 238894 435978
rect 238962 435922 239018 435978
rect 269558 436294 269614 436350
rect 269682 436294 269738 436350
rect 269558 436170 269614 436226
rect 269682 436170 269738 436226
rect 269558 436046 269614 436102
rect 269682 436046 269738 436102
rect 269558 435922 269614 435978
rect 269682 435922 269738 435978
rect 300278 436294 300334 436350
rect 300402 436294 300458 436350
rect 300278 436170 300334 436226
rect 300402 436170 300458 436226
rect 300278 436046 300334 436102
rect 300402 436046 300458 436102
rect 300278 435922 300334 435978
rect 300402 435922 300458 435978
rect 330998 436294 331054 436350
rect 331122 436294 331178 436350
rect 330998 436170 331054 436226
rect 331122 436170 331178 436226
rect 330998 436046 331054 436102
rect 331122 436046 331178 436102
rect 330998 435922 331054 435978
rect 331122 435922 331178 435978
rect 361718 436294 361774 436350
rect 361842 436294 361898 436350
rect 361718 436170 361774 436226
rect 361842 436170 361898 436226
rect 361718 436046 361774 436102
rect 361842 436046 361898 436102
rect 361718 435922 361774 435978
rect 361842 435922 361898 435978
rect 392438 436294 392494 436350
rect 392562 436294 392618 436350
rect 392438 436170 392494 436226
rect 392562 436170 392618 436226
rect 392438 436046 392494 436102
rect 392562 436046 392618 436102
rect 392438 435922 392494 435978
rect 392562 435922 392618 435978
rect 423158 436294 423214 436350
rect 423282 436294 423338 436350
rect 423158 436170 423214 436226
rect 423282 436170 423338 436226
rect 423158 436046 423214 436102
rect 423282 436046 423338 436102
rect 423158 435922 423214 435978
rect 423282 435922 423338 435978
rect 453878 436294 453934 436350
rect 454002 436294 454058 436350
rect 453878 436170 453934 436226
rect 454002 436170 454058 436226
rect 453878 436046 453934 436102
rect 454002 436046 454058 436102
rect 453878 435922 453934 435978
rect 454002 435922 454058 435978
rect 484598 436294 484654 436350
rect 484722 436294 484778 436350
rect 484598 436170 484654 436226
rect 484722 436170 484778 436226
rect 484598 436046 484654 436102
rect 484722 436046 484778 436102
rect 484598 435922 484654 435978
rect 484722 435922 484778 435978
rect 515318 436294 515374 436350
rect 515442 436294 515498 436350
rect 515318 436170 515374 436226
rect 515442 436170 515498 436226
rect 515318 436046 515374 436102
rect 515442 436046 515498 436102
rect 515318 435922 515374 435978
rect 515442 435922 515498 435978
rect 546038 436294 546094 436350
rect 546162 436294 546218 436350
rect 546038 436170 546094 436226
rect 546162 436170 546218 436226
rect 546038 436046 546094 436102
rect 546162 436046 546218 436102
rect 546038 435922 546094 435978
rect 546162 435922 546218 435978
rect 561250 436294 561306 436350
rect 561374 436294 561430 436350
rect 561498 436294 561554 436350
rect 561622 436294 561678 436350
rect 561250 436170 561306 436226
rect 561374 436170 561430 436226
rect 561498 436170 561554 436226
rect 561622 436170 561678 436226
rect 561250 436046 561306 436102
rect 561374 436046 561430 436102
rect 561498 436046 561554 436102
rect 561622 436046 561678 436102
rect 561250 435922 561306 435978
rect 561374 435922 561430 435978
rect 561498 435922 561554 435978
rect 561622 435922 561678 435978
rect 131318 424294 131374 424350
rect 131442 424294 131498 424350
rect 131318 424170 131374 424226
rect 131442 424170 131498 424226
rect 131318 424046 131374 424102
rect 131442 424046 131498 424102
rect 131318 423922 131374 423978
rect 131442 423922 131498 423978
rect 162038 424294 162094 424350
rect 162162 424294 162218 424350
rect 162038 424170 162094 424226
rect 162162 424170 162218 424226
rect 162038 424046 162094 424102
rect 162162 424046 162218 424102
rect 162038 423922 162094 423978
rect 162162 423922 162218 423978
rect 192758 424294 192814 424350
rect 192882 424294 192938 424350
rect 192758 424170 192814 424226
rect 192882 424170 192938 424226
rect 192758 424046 192814 424102
rect 192882 424046 192938 424102
rect 192758 423922 192814 423978
rect 192882 423922 192938 423978
rect 223478 424294 223534 424350
rect 223602 424294 223658 424350
rect 223478 424170 223534 424226
rect 223602 424170 223658 424226
rect 223478 424046 223534 424102
rect 223602 424046 223658 424102
rect 223478 423922 223534 423978
rect 223602 423922 223658 423978
rect 254198 424294 254254 424350
rect 254322 424294 254378 424350
rect 254198 424170 254254 424226
rect 254322 424170 254378 424226
rect 254198 424046 254254 424102
rect 254322 424046 254378 424102
rect 254198 423922 254254 423978
rect 254322 423922 254378 423978
rect 284918 424294 284974 424350
rect 285042 424294 285098 424350
rect 284918 424170 284974 424226
rect 285042 424170 285098 424226
rect 284918 424046 284974 424102
rect 285042 424046 285098 424102
rect 284918 423922 284974 423978
rect 285042 423922 285098 423978
rect 315638 424294 315694 424350
rect 315762 424294 315818 424350
rect 315638 424170 315694 424226
rect 315762 424170 315818 424226
rect 315638 424046 315694 424102
rect 315762 424046 315818 424102
rect 315638 423922 315694 423978
rect 315762 423922 315818 423978
rect 346358 424294 346414 424350
rect 346482 424294 346538 424350
rect 346358 424170 346414 424226
rect 346482 424170 346538 424226
rect 346358 424046 346414 424102
rect 346482 424046 346538 424102
rect 346358 423922 346414 423978
rect 346482 423922 346538 423978
rect 377078 424294 377134 424350
rect 377202 424294 377258 424350
rect 377078 424170 377134 424226
rect 377202 424170 377258 424226
rect 377078 424046 377134 424102
rect 377202 424046 377258 424102
rect 377078 423922 377134 423978
rect 377202 423922 377258 423978
rect 407798 424294 407854 424350
rect 407922 424294 407978 424350
rect 407798 424170 407854 424226
rect 407922 424170 407978 424226
rect 407798 424046 407854 424102
rect 407922 424046 407978 424102
rect 407798 423922 407854 423978
rect 407922 423922 407978 423978
rect 438518 424294 438574 424350
rect 438642 424294 438698 424350
rect 438518 424170 438574 424226
rect 438642 424170 438698 424226
rect 438518 424046 438574 424102
rect 438642 424046 438698 424102
rect 438518 423922 438574 423978
rect 438642 423922 438698 423978
rect 469238 424294 469294 424350
rect 469362 424294 469418 424350
rect 469238 424170 469294 424226
rect 469362 424170 469418 424226
rect 469238 424046 469294 424102
rect 469362 424046 469418 424102
rect 469238 423922 469294 423978
rect 469362 423922 469418 423978
rect 499958 424294 500014 424350
rect 500082 424294 500138 424350
rect 499958 424170 500014 424226
rect 500082 424170 500138 424226
rect 499958 424046 500014 424102
rect 500082 424046 500138 424102
rect 499958 423922 500014 423978
rect 500082 423922 500138 423978
rect 530678 424294 530734 424350
rect 530802 424294 530858 424350
rect 530678 424170 530734 424226
rect 530802 424170 530858 424226
rect 530678 424046 530734 424102
rect 530802 424046 530858 424102
rect 530678 423922 530734 423978
rect 530802 423922 530858 423978
rect 111250 418294 111306 418350
rect 111374 418294 111430 418350
rect 111498 418294 111554 418350
rect 111622 418294 111678 418350
rect 111250 418170 111306 418226
rect 111374 418170 111430 418226
rect 111498 418170 111554 418226
rect 111622 418170 111678 418226
rect 111250 418046 111306 418102
rect 111374 418046 111430 418102
rect 111498 418046 111554 418102
rect 111622 418046 111678 418102
rect 111250 417922 111306 417978
rect 111374 417922 111430 417978
rect 111498 417922 111554 417978
rect 111622 417922 111678 417978
rect 96970 406294 97026 406350
rect 97094 406294 97150 406350
rect 97218 406294 97274 406350
rect 97342 406294 97398 406350
rect 96970 406170 97026 406226
rect 97094 406170 97150 406226
rect 97218 406170 97274 406226
rect 97342 406170 97398 406226
rect 96970 406046 97026 406102
rect 97094 406046 97150 406102
rect 97218 406046 97274 406102
rect 97342 406046 97398 406102
rect 96970 405922 97026 405978
rect 97094 405922 97150 405978
rect 97218 405922 97274 405978
rect 97342 405922 97398 405978
rect 100598 406294 100654 406350
rect 100722 406294 100778 406350
rect 100598 406170 100654 406226
rect 100722 406170 100778 406226
rect 100598 406046 100654 406102
rect 100722 406046 100778 406102
rect 100598 405922 100654 405978
rect 100722 405922 100778 405978
rect 115958 418294 116014 418350
rect 116082 418294 116138 418350
rect 115958 418170 116014 418226
rect 116082 418170 116138 418226
rect 115958 418046 116014 418102
rect 116082 418046 116138 418102
rect 115958 417922 116014 417978
rect 116082 417922 116138 417978
rect 146678 418294 146734 418350
rect 146802 418294 146858 418350
rect 146678 418170 146734 418226
rect 146802 418170 146858 418226
rect 146678 418046 146734 418102
rect 146802 418046 146858 418102
rect 146678 417922 146734 417978
rect 146802 417922 146858 417978
rect 177398 418294 177454 418350
rect 177522 418294 177578 418350
rect 177398 418170 177454 418226
rect 177522 418170 177578 418226
rect 177398 418046 177454 418102
rect 177522 418046 177578 418102
rect 177398 417922 177454 417978
rect 177522 417922 177578 417978
rect 208118 418294 208174 418350
rect 208242 418294 208298 418350
rect 208118 418170 208174 418226
rect 208242 418170 208298 418226
rect 208118 418046 208174 418102
rect 208242 418046 208298 418102
rect 208118 417922 208174 417978
rect 208242 417922 208298 417978
rect 238838 418294 238894 418350
rect 238962 418294 239018 418350
rect 238838 418170 238894 418226
rect 238962 418170 239018 418226
rect 238838 418046 238894 418102
rect 238962 418046 239018 418102
rect 238838 417922 238894 417978
rect 238962 417922 239018 417978
rect 269558 418294 269614 418350
rect 269682 418294 269738 418350
rect 269558 418170 269614 418226
rect 269682 418170 269738 418226
rect 269558 418046 269614 418102
rect 269682 418046 269738 418102
rect 269558 417922 269614 417978
rect 269682 417922 269738 417978
rect 300278 418294 300334 418350
rect 300402 418294 300458 418350
rect 300278 418170 300334 418226
rect 300402 418170 300458 418226
rect 300278 418046 300334 418102
rect 300402 418046 300458 418102
rect 300278 417922 300334 417978
rect 300402 417922 300458 417978
rect 330998 418294 331054 418350
rect 331122 418294 331178 418350
rect 330998 418170 331054 418226
rect 331122 418170 331178 418226
rect 330998 418046 331054 418102
rect 331122 418046 331178 418102
rect 330998 417922 331054 417978
rect 331122 417922 331178 417978
rect 361718 418294 361774 418350
rect 361842 418294 361898 418350
rect 361718 418170 361774 418226
rect 361842 418170 361898 418226
rect 361718 418046 361774 418102
rect 361842 418046 361898 418102
rect 361718 417922 361774 417978
rect 361842 417922 361898 417978
rect 392438 418294 392494 418350
rect 392562 418294 392618 418350
rect 392438 418170 392494 418226
rect 392562 418170 392618 418226
rect 392438 418046 392494 418102
rect 392562 418046 392618 418102
rect 392438 417922 392494 417978
rect 392562 417922 392618 417978
rect 423158 418294 423214 418350
rect 423282 418294 423338 418350
rect 423158 418170 423214 418226
rect 423282 418170 423338 418226
rect 423158 418046 423214 418102
rect 423282 418046 423338 418102
rect 423158 417922 423214 417978
rect 423282 417922 423338 417978
rect 453878 418294 453934 418350
rect 454002 418294 454058 418350
rect 453878 418170 453934 418226
rect 454002 418170 454058 418226
rect 453878 418046 453934 418102
rect 454002 418046 454058 418102
rect 453878 417922 453934 417978
rect 454002 417922 454058 417978
rect 484598 418294 484654 418350
rect 484722 418294 484778 418350
rect 484598 418170 484654 418226
rect 484722 418170 484778 418226
rect 484598 418046 484654 418102
rect 484722 418046 484778 418102
rect 484598 417922 484654 417978
rect 484722 417922 484778 417978
rect 515318 418294 515374 418350
rect 515442 418294 515498 418350
rect 515318 418170 515374 418226
rect 515442 418170 515498 418226
rect 515318 418046 515374 418102
rect 515442 418046 515498 418102
rect 515318 417922 515374 417978
rect 515442 417922 515498 417978
rect 546038 418294 546094 418350
rect 546162 418294 546218 418350
rect 546038 418170 546094 418226
rect 546162 418170 546218 418226
rect 546038 418046 546094 418102
rect 546162 418046 546218 418102
rect 546038 417922 546094 417978
rect 546162 417922 546218 417978
rect 561250 418294 561306 418350
rect 561374 418294 561430 418350
rect 561498 418294 561554 418350
rect 561622 418294 561678 418350
rect 561250 418170 561306 418226
rect 561374 418170 561430 418226
rect 561498 418170 561554 418226
rect 561622 418170 561678 418226
rect 561250 418046 561306 418102
rect 561374 418046 561430 418102
rect 561498 418046 561554 418102
rect 561622 418046 561678 418102
rect 561250 417922 561306 417978
rect 561374 417922 561430 417978
rect 561498 417922 561554 417978
rect 561622 417922 561678 417978
rect 131318 406294 131374 406350
rect 131442 406294 131498 406350
rect 131318 406170 131374 406226
rect 131442 406170 131498 406226
rect 131318 406046 131374 406102
rect 131442 406046 131498 406102
rect 131318 405922 131374 405978
rect 131442 405922 131498 405978
rect 162038 406294 162094 406350
rect 162162 406294 162218 406350
rect 162038 406170 162094 406226
rect 162162 406170 162218 406226
rect 162038 406046 162094 406102
rect 162162 406046 162218 406102
rect 162038 405922 162094 405978
rect 162162 405922 162218 405978
rect 192758 406294 192814 406350
rect 192882 406294 192938 406350
rect 192758 406170 192814 406226
rect 192882 406170 192938 406226
rect 192758 406046 192814 406102
rect 192882 406046 192938 406102
rect 192758 405922 192814 405978
rect 192882 405922 192938 405978
rect 223478 406294 223534 406350
rect 223602 406294 223658 406350
rect 223478 406170 223534 406226
rect 223602 406170 223658 406226
rect 223478 406046 223534 406102
rect 223602 406046 223658 406102
rect 223478 405922 223534 405978
rect 223602 405922 223658 405978
rect 254198 406294 254254 406350
rect 254322 406294 254378 406350
rect 254198 406170 254254 406226
rect 254322 406170 254378 406226
rect 254198 406046 254254 406102
rect 254322 406046 254378 406102
rect 254198 405922 254254 405978
rect 254322 405922 254378 405978
rect 284918 406294 284974 406350
rect 285042 406294 285098 406350
rect 284918 406170 284974 406226
rect 285042 406170 285098 406226
rect 284918 406046 284974 406102
rect 285042 406046 285098 406102
rect 284918 405922 284974 405978
rect 285042 405922 285098 405978
rect 315638 406294 315694 406350
rect 315762 406294 315818 406350
rect 315638 406170 315694 406226
rect 315762 406170 315818 406226
rect 315638 406046 315694 406102
rect 315762 406046 315818 406102
rect 315638 405922 315694 405978
rect 315762 405922 315818 405978
rect 346358 406294 346414 406350
rect 346482 406294 346538 406350
rect 346358 406170 346414 406226
rect 346482 406170 346538 406226
rect 346358 406046 346414 406102
rect 346482 406046 346538 406102
rect 346358 405922 346414 405978
rect 346482 405922 346538 405978
rect 377078 406294 377134 406350
rect 377202 406294 377258 406350
rect 377078 406170 377134 406226
rect 377202 406170 377258 406226
rect 377078 406046 377134 406102
rect 377202 406046 377258 406102
rect 377078 405922 377134 405978
rect 377202 405922 377258 405978
rect 407798 406294 407854 406350
rect 407922 406294 407978 406350
rect 407798 406170 407854 406226
rect 407922 406170 407978 406226
rect 407798 406046 407854 406102
rect 407922 406046 407978 406102
rect 407798 405922 407854 405978
rect 407922 405922 407978 405978
rect 438518 406294 438574 406350
rect 438642 406294 438698 406350
rect 438518 406170 438574 406226
rect 438642 406170 438698 406226
rect 438518 406046 438574 406102
rect 438642 406046 438698 406102
rect 438518 405922 438574 405978
rect 438642 405922 438698 405978
rect 469238 406294 469294 406350
rect 469362 406294 469418 406350
rect 469238 406170 469294 406226
rect 469362 406170 469418 406226
rect 469238 406046 469294 406102
rect 469362 406046 469418 406102
rect 469238 405922 469294 405978
rect 469362 405922 469418 405978
rect 499958 406294 500014 406350
rect 500082 406294 500138 406350
rect 499958 406170 500014 406226
rect 500082 406170 500138 406226
rect 499958 406046 500014 406102
rect 500082 406046 500138 406102
rect 499958 405922 500014 405978
rect 500082 405922 500138 405978
rect 530678 406294 530734 406350
rect 530802 406294 530858 406350
rect 530678 406170 530734 406226
rect 530802 406170 530858 406226
rect 530678 406046 530734 406102
rect 530802 406046 530858 406102
rect 530678 405922 530734 405978
rect 530802 405922 530858 405978
rect 111250 400294 111306 400350
rect 111374 400294 111430 400350
rect 111498 400294 111554 400350
rect 111622 400294 111678 400350
rect 111250 400170 111306 400226
rect 111374 400170 111430 400226
rect 111498 400170 111554 400226
rect 111622 400170 111678 400226
rect 111250 400046 111306 400102
rect 111374 400046 111430 400102
rect 111498 400046 111554 400102
rect 111622 400046 111678 400102
rect 111250 399922 111306 399978
rect 111374 399922 111430 399978
rect 111498 399922 111554 399978
rect 111622 399922 111678 399978
rect 96970 388294 97026 388350
rect 97094 388294 97150 388350
rect 97218 388294 97274 388350
rect 97342 388294 97398 388350
rect 96970 388170 97026 388226
rect 97094 388170 97150 388226
rect 97218 388170 97274 388226
rect 97342 388170 97398 388226
rect 96970 388046 97026 388102
rect 97094 388046 97150 388102
rect 97218 388046 97274 388102
rect 97342 388046 97398 388102
rect 96970 387922 97026 387978
rect 97094 387922 97150 387978
rect 97218 387922 97274 387978
rect 97342 387922 97398 387978
rect 100598 388294 100654 388350
rect 100722 388294 100778 388350
rect 100598 388170 100654 388226
rect 100722 388170 100778 388226
rect 100598 388046 100654 388102
rect 100722 388046 100778 388102
rect 100598 387922 100654 387978
rect 100722 387922 100778 387978
rect 115958 400294 116014 400350
rect 116082 400294 116138 400350
rect 115958 400170 116014 400226
rect 116082 400170 116138 400226
rect 115958 400046 116014 400102
rect 116082 400046 116138 400102
rect 115958 399922 116014 399978
rect 116082 399922 116138 399978
rect 146678 400294 146734 400350
rect 146802 400294 146858 400350
rect 146678 400170 146734 400226
rect 146802 400170 146858 400226
rect 146678 400046 146734 400102
rect 146802 400046 146858 400102
rect 146678 399922 146734 399978
rect 146802 399922 146858 399978
rect 177398 400294 177454 400350
rect 177522 400294 177578 400350
rect 177398 400170 177454 400226
rect 177522 400170 177578 400226
rect 177398 400046 177454 400102
rect 177522 400046 177578 400102
rect 177398 399922 177454 399978
rect 177522 399922 177578 399978
rect 208118 400294 208174 400350
rect 208242 400294 208298 400350
rect 208118 400170 208174 400226
rect 208242 400170 208298 400226
rect 208118 400046 208174 400102
rect 208242 400046 208298 400102
rect 208118 399922 208174 399978
rect 208242 399922 208298 399978
rect 238838 400294 238894 400350
rect 238962 400294 239018 400350
rect 238838 400170 238894 400226
rect 238962 400170 239018 400226
rect 238838 400046 238894 400102
rect 238962 400046 239018 400102
rect 238838 399922 238894 399978
rect 238962 399922 239018 399978
rect 269558 400294 269614 400350
rect 269682 400294 269738 400350
rect 269558 400170 269614 400226
rect 269682 400170 269738 400226
rect 269558 400046 269614 400102
rect 269682 400046 269738 400102
rect 269558 399922 269614 399978
rect 269682 399922 269738 399978
rect 300278 400294 300334 400350
rect 300402 400294 300458 400350
rect 300278 400170 300334 400226
rect 300402 400170 300458 400226
rect 300278 400046 300334 400102
rect 300402 400046 300458 400102
rect 300278 399922 300334 399978
rect 300402 399922 300458 399978
rect 330998 400294 331054 400350
rect 331122 400294 331178 400350
rect 330998 400170 331054 400226
rect 331122 400170 331178 400226
rect 330998 400046 331054 400102
rect 331122 400046 331178 400102
rect 330998 399922 331054 399978
rect 331122 399922 331178 399978
rect 361718 400294 361774 400350
rect 361842 400294 361898 400350
rect 361718 400170 361774 400226
rect 361842 400170 361898 400226
rect 361718 400046 361774 400102
rect 361842 400046 361898 400102
rect 361718 399922 361774 399978
rect 361842 399922 361898 399978
rect 392438 400294 392494 400350
rect 392562 400294 392618 400350
rect 392438 400170 392494 400226
rect 392562 400170 392618 400226
rect 392438 400046 392494 400102
rect 392562 400046 392618 400102
rect 392438 399922 392494 399978
rect 392562 399922 392618 399978
rect 423158 400294 423214 400350
rect 423282 400294 423338 400350
rect 423158 400170 423214 400226
rect 423282 400170 423338 400226
rect 423158 400046 423214 400102
rect 423282 400046 423338 400102
rect 423158 399922 423214 399978
rect 423282 399922 423338 399978
rect 453878 400294 453934 400350
rect 454002 400294 454058 400350
rect 453878 400170 453934 400226
rect 454002 400170 454058 400226
rect 453878 400046 453934 400102
rect 454002 400046 454058 400102
rect 453878 399922 453934 399978
rect 454002 399922 454058 399978
rect 484598 400294 484654 400350
rect 484722 400294 484778 400350
rect 484598 400170 484654 400226
rect 484722 400170 484778 400226
rect 484598 400046 484654 400102
rect 484722 400046 484778 400102
rect 484598 399922 484654 399978
rect 484722 399922 484778 399978
rect 515318 400294 515374 400350
rect 515442 400294 515498 400350
rect 515318 400170 515374 400226
rect 515442 400170 515498 400226
rect 515318 400046 515374 400102
rect 515442 400046 515498 400102
rect 515318 399922 515374 399978
rect 515442 399922 515498 399978
rect 546038 400294 546094 400350
rect 546162 400294 546218 400350
rect 546038 400170 546094 400226
rect 546162 400170 546218 400226
rect 546038 400046 546094 400102
rect 546162 400046 546218 400102
rect 546038 399922 546094 399978
rect 546162 399922 546218 399978
rect 561250 400294 561306 400350
rect 561374 400294 561430 400350
rect 561498 400294 561554 400350
rect 561622 400294 561678 400350
rect 561250 400170 561306 400226
rect 561374 400170 561430 400226
rect 561498 400170 561554 400226
rect 561622 400170 561678 400226
rect 561250 400046 561306 400102
rect 561374 400046 561430 400102
rect 561498 400046 561554 400102
rect 561622 400046 561678 400102
rect 561250 399922 561306 399978
rect 561374 399922 561430 399978
rect 561498 399922 561554 399978
rect 561622 399922 561678 399978
rect 131318 388294 131374 388350
rect 131442 388294 131498 388350
rect 131318 388170 131374 388226
rect 131442 388170 131498 388226
rect 131318 388046 131374 388102
rect 131442 388046 131498 388102
rect 131318 387922 131374 387978
rect 131442 387922 131498 387978
rect 162038 388294 162094 388350
rect 162162 388294 162218 388350
rect 162038 388170 162094 388226
rect 162162 388170 162218 388226
rect 162038 388046 162094 388102
rect 162162 388046 162218 388102
rect 162038 387922 162094 387978
rect 162162 387922 162218 387978
rect 192758 388294 192814 388350
rect 192882 388294 192938 388350
rect 192758 388170 192814 388226
rect 192882 388170 192938 388226
rect 192758 388046 192814 388102
rect 192882 388046 192938 388102
rect 192758 387922 192814 387978
rect 192882 387922 192938 387978
rect 223478 388294 223534 388350
rect 223602 388294 223658 388350
rect 223478 388170 223534 388226
rect 223602 388170 223658 388226
rect 223478 388046 223534 388102
rect 223602 388046 223658 388102
rect 223478 387922 223534 387978
rect 223602 387922 223658 387978
rect 254198 388294 254254 388350
rect 254322 388294 254378 388350
rect 254198 388170 254254 388226
rect 254322 388170 254378 388226
rect 254198 388046 254254 388102
rect 254322 388046 254378 388102
rect 254198 387922 254254 387978
rect 254322 387922 254378 387978
rect 284918 388294 284974 388350
rect 285042 388294 285098 388350
rect 284918 388170 284974 388226
rect 285042 388170 285098 388226
rect 284918 388046 284974 388102
rect 285042 388046 285098 388102
rect 284918 387922 284974 387978
rect 285042 387922 285098 387978
rect 315638 388294 315694 388350
rect 315762 388294 315818 388350
rect 315638 388170 315694 388226
rect 315762 388170 315818 388226
rect 315638 388046 315694 388102
rect 315762 388046 315818 388102
rect 315638 387922 315694 387978
rect 315762 387922 315818 387978
rect 346358 388294 346414 388350
rect 346482 388294 346538 388350
rect 346358 388170 346414 388226
rect 346482 388170 346538 388226
rect 346358 388046 346414 388102
rect 346482 388046 346538 388102
rect 346358 387922 346414 387978
rect 346482 387922 346538 387978
rect 377078 388294 377134 388350
rect 377202 388294 377258 388350
rect 377078 388170 377134 388226
rect 377202 388170 377258 388226
rect 377078 388046 377134 388102
rect 377202 388046 377258 388102
rect 377078 387922 377134 387978
rect 377202 387922 377258 387978
rect 407798 388294 407854 388350
rect 407922 388294 407978 388350
rect 407798 388170 407854 388226
rect 407922 388170 407978 388226
rect 407798 388046 407854 388102
rect 407922 388046 407978 388102
rect 407798 387922 407854 387978
rect 407922 387922 407978 387978
rect 438518 388294 438574 388350
rect 438642 388294 438698 388350
rect 438518 388170 438574 388226
rect 438642 388170 438698 388226
rect 438518 388046 438574 388102
rect 438642 388046 438698 388102
rect 438518 387922 438574 387978
rect 438642 387922 438698 387978
rect 469238 388294 469294 388350
rect 469362 388294 469418 388350
rect 469238 388170 469294 388226
rect 469362 388170 469418 388226
rect 469238 388046 469294 388102
rect 469362 388046 469418 388102
rect 469238 387922 469294 387978
rect 469362 387922 469418 387978
rect 499958 388294 500014 388350
rect 500082 388294 500138 388350
rect 499958 388170 500014 388226
rect 500082 388170 500138 388226
rect 499958 388046 500014 388102
rect 500082 388046 500138 388102
rect 499958 387922 500014 387978
rect 500082 387922 500138 387978
rect 530678 388294 530734 388350
rect 530802 388294 530858 388350
rect 530678 388170 530734 388226
rect 530802 388170 530858 388226
rect 530678 388046 530734 388102
rect 530802 388046 530858 388102
rect 530678 387922 530734 387978
rect 530802 387922 530858 387978
rect 111250 382294 111306 382350
rect 111374 382294 111430 382350
rect 111498 382294 111554 382350
rect 111622 382294 111678 382350
rect 111250 382170 111306 382226
rect 111374 382170 111430 382226
rect 111498 382170 111554 382226
rect 111622 382170 111678 382226
rect 111250 382046 111306 382102
rect 111374 382046 111430 382102
rect 111498 382046 111554 382102
rect 111622 382046 111678 382102
rect 111250 381922 111306 381978
rect 111374 381922 111430 381978
rect 111498 381922 111554 381978
rect 111622 381922 111678 381978
rect 96970 370294 97026 370350
rect 97094 370294 97150 370350
rect 97218 370294 97274 370350
rect 97342 370294 97398 370350
rect 96970 370170 97026 370226
rect 97094 370170 97150 370226
rect 97218 370170 97274 370226
rect 97342 370170 97398 370226
rect 96970 370046 97026 370102
rect 97094 370046 97150 370102
rect 97218 370046 97274 370102
rect 97342 370046 97398 370102
rect 96970 369922 97026 369978
rect 97094 369922 97150 369978
rect 97218 369922 97274 369978
rect 97342 369922 97398 369978
rect 100598 370294 100654 370350
rect 100722 370294 100778 370350
rect 100598 370170 100654 370226
rect 100722 370170 100778 370226
rect 100598 370046 100654 370102
rect 100722 370046 100778 370102
rect 100598 369922 100654 369978
rect 100722 369922 100778 369978
rect 115958 382294 116014 382350
rect 116082 382294 116138 382350
rect 115958 382170 116014 382226
rect 116082 382170 116138 382226
rect 115958 382046 116014 382102
rect 116082 382046 116138 382102
rect 115958 381922 116014 381978
rect 116082 381922 116138 381978
rect 146678 382294 146734 382350
rect 146802 382294 146858 382350
rect 146678 382170 146734 382226
rect 146802 382170 146858 382226
rect 146678 382046 146734 382102
rect 146802 382046 146858 382102
rect 146678 381922 146734 381978
rect 146802 381922 146858 381978
rect 177398 382294 177454 382350
rect 177522 382294 177578 382350
rect 177398 382170 177454 382226
rect 177522 382170 177578 382226
rect 177398 382046 177454 382102
rect 177522 382046 177578 382102
rect 177398 381922 177454 381978
rect 177522 381922 177578 381978
rect 208118 382294 208174 382350
rect 208242 382294 208298 382350
rect 208118 382170 208174 382226
rect 208242 382170 208298 382226
rect 208118 382046 208174 382102
rect 208242 382046 208298 382102
rect 208118 381922 208174 381978
rect 208242 381922 208298 381978
rect 238838 382294 238894 382350
rect 238962 382294 239018 382350
rect 238838 382170 238894 382226
rect 238962 382170 239018 382226
rect 238838 382046 238894 382102
rect 238962 382046 239018 382102
rect 238838 381922 238894 381978
rect 238962 381922 239018 381978
rect 269558 382294 269614 382350
rect 269682 382294 269738 382350
rect 269558 382170 269614 382226
rect 269682 382170 269738 382226
rect 269558 382046 269614 382102
rect 269682 382046 269738 382102
rect 269558 381922 269614 381978
rect 269682 381922 269738 381978
rect 300278 382294 300334 382350
rect 300402 382294 300458 382350
rect 300278 382170 300334 382226
rect 300402 382170 300458 382226
rect 300278 382046 300334 382102
rect 300402 382046 300458 382102
rect 300278 381922 300334 381978
rect 300402 381922 300458 381978
rect 330998 382294 331054 382350
rect 331122 382294 331178 382350
rect 330998 382170 331054 382226
rect 331122 382170 331178 382226
rect 330998 382046 331054 382102
rect 331122 382046 331178 382102
rect 330998 381922 331054 381978
rect 331122 381922 331178 381978
rect 361718 382294 361774 382350
rect 361842 382294 361898 382350
rect 361718 382170 361774 382226
rect 361842 382170 361898 382226
rect 361718 382046 361774 382102
rect 361842 382046 361898 382102
rect 361718 381922 361774 381978
rect 361842 381922 361898 381978
rect 392438 382294 392494 382350
rect 392562 382294 392618 382350
rect 392438 382170 392494 382226
rect 392562 382170 392618 382226
rect 392438 382046 392494 382102
rect 392562 382046 392618 382102
rect 392438 381922 392494 381978
rect 392562 381922 392618 381978
rect 423158 382294 423214 382350
rect 423282 382294 423338 382350
rect 423158 382170 423214 382226
rect 423282 382170 423338 382226
rect 423158 382046 423214 382102
rect 423282 382046 423338 382102
rect 423158 381922 423214 381978
rect 423282 381922 423338 381978
rect 453878 382294 453934 382350
rect 454002 382294 454058 382350
rect 453878 382170 453934 382226
rect 454002 382170 454058 382226
rect 453878 382046 453934 382102
rect 454002 382046 454058 382102
rect 453878 381922 453934 381978
rect 454002 381922 454058 381978
rect 484598 382294 484654 382350
rect 484722 382294 484778 382350
rect 484598 382170 484654 382226
rect 484722 382170 484778 382226
rect 484598 382046 484654 382102
rect 484722 382046 484778 382102
rect 484598 381922 484654 381978
rect 484722 381922 484778 381978
rect 515318 382294 515374 382350
rect 515442 382294 515498 382350
rect 515318 382170 515374 382226
rect 515442 382170 515498 382226
rect 515318 382046 515374 382102
rect 515442 382046 515498 382102
rect 515318 381922 515374 381978
rect 515442 381922 515498 381978
rect 546038 382294 546094 382350
rect 546162 382294 546218 382350
rect 546038 382170 546094 382226
rect 546162 382170 546218 382226
rect 546038 382046 546094 382102
rect 546162 382046 546218 382102
rect 546038 381922 546094 381978
rect 546162 381922 546218 381978
rect 561250 382294 561306 382350
rect 561374 382294 561430 382350
rect 561498 382294 561554 382350
rect 561622 382294 561678 382350
rect 561250 382170 561306 382226
rect 561374 382170 561430 382226
rect 561498 382170 561554 382226
rect 561622 382170 561678 382226
rect 561250 382046 561306 382102
rect 561374 382046 561430 382102
rect 561498 382046 561554 382102
rect 561622 382046 561678 382102
rect 561250 381922 561306 381978
rect 561374 381922 561430 381978
rect 561498 381922 561554 381978
rect 561622 381922 561678 381978
rect 131318 370294 131374 370350
rect 131442 370294 131498 370350
rect 131318 370170 131374 370226
rect 131442 370170 131498 370226
rect 131318 370046 131374 370102
rect 131442 370046 131498 370102
rect 131318 369922 131374 369978
rect 131442 369922 131498 369978
rect 162038 370294 162094 370350
rect 162162 370294 162218 370350
rect 162038 370170 162094 370226
rect 162162 370170 162218 370226
rect 162038 370046 162094 370102
rect 162162 370046 162218 370102
rect 162038 369922 162094 369978
rect 162162 369922 162218 369978
rect 192758 370294 192814 370350
rect 192882 370294 192938 370350
rect 192758 370170 192814 370226
rect 192882 370170 192938 370226
rect 192758 370046 192814 370102
rect 192882 370046 192938 370102
rect 192758 369922 192814 369978
rect 192882 369922 192938 369978
rect 223478 370294 223534 370350
rect 223602 370294 223658 370350
rect 223478 370170 223534 370226
rect 223602 370170 223658 370226
rect 223478 370046 223534 370102
rect 223602 370046 223658 370102
rect 223478 369922 223534 369978
rect 223602 369922 223658 369978
rect 254198 370294 254254 370350
rect 254322 370294 254378 370350
rect 254198 370170 254254 370226
rect 254322 370170 254378 370226
rect 254198 370046 254254 370102
rect 254322 370046 254378 370102
rect 254198 369922 254254 369978
rect 254322 369922 254378 369978
rect 284918 370294 284974 370350
rect 285042 370294 285098 370350
rect 284918 370170 284974 370226
rect 285042 370170 285098 370226
rect 284918 370046 284974 370102
rect 285042 370046 285098 370102
rect 284918 369922 284974 369978
rect 285042 369922 285098 369978
rect 315638 370294 315694 370350
rect 315762 370294 315818 370350
rect 315638 370170 315694 370226
rect 315762 370170 315818 370226
rect 315638 370046 315694 370102
rect 315762 370046 315818 370102
rect 315638 369922 315694 369978
rect 315762 369922 315818 369978
rect 346358 370294 346414 370350
rect 346482 370294 346538 370350
rect 346358 370170 346414 370226
rect 346482 370170 346538 370226
rect 346358 370046 346414 370102
rect 346482 370046 346538 370102
rect 346358 369922 346414 369978
rect 346482 369922 346538 369978
rect 377078 370294 377134 370350
rect 377202 370294 377258 370350
rect 377078 370170 377134 370226
rect 377202 370170 377258 370226
rect 377078 370046 377134 370102
rect 377202 370046 377258 370102
rect 377078 369922 377134 369978
rect 377202 369922 377258 369978
rect 407798 370294 407854 370350
rect 407922 370294 407978 370350
rect 407798 370170 407854 370226
rect 407922 370170 407978 370226
rect 407798 370046 407854 370102
rect 407922 370046 407978 370102
rect 407798 369922 407854 369978
rect 407922 369922 407978 369978
rect 438518 370294 438574 370350
rect 438642 370294 438698 370350
rect 438518 370170 438574 370226
rect 438642 370170 438698 370226
rect 438518 370046 438574 370102
rect 438642 370046 438698 370102
rect 438518 369922 438574 369978
rect 438642 369922 438698 369978
rect 469238 370294 469294 370350
rect 469362 370294 469418 370350
rect 469238 370170 469294 370226
rect 469362 370170 469418 370226
rect 469238 370046 469294 370102
rect 469362 370046 469418 370102
rect 469238 369922 469294 369978
rect 469362 369922 469418 369978
rect 499958 370294 500014 370350
rect 500082 370294 500138 370350
rect 499958 370170 500014 370226
rect 500082 370170 500138 370226
rect 499958 370046 500014 370102
rect 500082 370046 500138 370102
rect 499958 369922 500014 369978
rect 500082 369922 500138 369978
rect 530678 370294 530734 370350
rect 530802 370294 530858 370350
rect 530678 370170 530734 370226
rect 530802 370170 530858 370226
rect 530678 370046 530734 370102
rect 530802 370046 530858 370102
rect 530678 369922 530734 369978
rect 530802 369922 530858 369978
rect 111250 364294 111306 364350
rect 111374 364294 111430 364350
rect 111498 364294 111554 364350
rect 111622 364294 111678 364350
rect 111250 364170 111306 364226
rect 111374 364170 111430 364226
rect 111498 364170 111554 364226
rect 111622 364170 111678 364226
rect 111250 364046 111306 364102
rect 111374 364046 111430 364102
rect 111498 364046 111554 364102
rect 111622 364046 111678 364102
rect 111250 363922 111306 363978
rect 111374 363922 111430 363978
rect 111498 363922 111554 363978
rect 111622 363922 111678 363978
rect 96970 352294 97026 352350
rect 97094 352294 97150 352350
rect 97218 352294 97274 352350
rect 97342 352294 97398 352350
rect 96970 352170 97026 352226
rect 97094 352170 97150 352226
rect 97218 352170 97274 352226
rect 97342 352170 97398 352226
rect 96970 352046 97026 352102
rect 97094 352046 97150 352102
rect 97218 352046 97274 352102
rect 97342 352046 97398 352102
rect 96970 351922 97026 351978
rect 97094 351922 97150 351978
rect 97218 351922 97274 351978
rect 97342 351922 97398 351978
rect 100598 352294 100654 352350
rect 100722 352294 100778 352350
rect 100598 352170 100654 352226
rect 100722 352170 100778 352226
rect 100598 352046 100654 352102
rect 100722 352046 100778 352102
rect 100598 351922 100654 351978
rect 100722 351922 100778 351978
rect 115958 364294 116014 364350
rect 116082 364294 116138 364350
rect 115958 364170 116014 364226
rect 116082 364170 116138 364226
rect 115958 364046 116014 364102
rect 116082 364046 116138 364102
rect 115958 363922 116014 363978
rect 116082 363922 116138 363978
rect 146678 364294 146734 364350
rect 146802 364294 146858 364350
rect 146678 364170 146734 364226
rect 146802 364170 146858 364226
rect 146678 364046 146734 364102
rect 146802 364046 146858 364102
rect 146678 363922 146734 363978
rect 146802 363922 146858 363978
rect 177398 364294 177454 364350
rect 177522 364294 177578 364350
rect 177398 364170 177454 364226
rect 177522 364170 177578 364226
rect 177398 364046 177454 364102
rect 177522 364046 177578 364102
rect 177398 363922 177454 363978
rect 177522 363922 177578 363978
rect 208118 364294 208174 364350
rect 208242 364294 208298 364350
rect 208118 364170 208174 364226
rect 208242 364170 208298 364226
rect 208118 364046 208174 364102
rect 208242 364046 208298 364102
rect 208118 363922 208174 363978
rect 208242 363922 208298 363978
rect 238838 364294 238894 364350
rect 238962 364294 239018 364350
rect 238838 364170 238894 364226
rect 238962 364170 239018 364226
rect 238838 364046 238894 364102
rect 238962 364046 239018 364102
rect 238838 363922 238894 363978
rect 238962 363922 239018 363978
rect 269558 364294 269614 364350
rect 269682 364294 269738 364350
rect 269558 364170 269614 364226
rect 269682 364170 269738 364226
rect 269558 364046 269614 364102
rect 269682 364046 269738 364102
rect 269558 363922 269614 363978
rect 269682 363922 269738 363978
rect 300278 364294 300334 364350
rect 300402 364294 300458 364350
rect 300278 364170 300334 364226
rect 300402 364170 300458 364226
rect 300278 364046 300334 364102
rect 300402 364046 300458 364102
rect 300278 363922 300334 363978
rect 300402 363922 300458 363978
rect 330998 364294 331054 364350
rect 331122 364294 331178 364350
rect 330998 364170 331054 364226
rect 331122 364170 331178 364226
rect 330998 364046 331054 364102
rect 331122 364046 331178 364102
rect 330998 363922 331054 363978
rect 331122 363922 331178 363978
rect 361718 364294 361774 364350
rect 361842 364294 361898 364350
rect 361718 364170 361774 364226
rect 361842 364170 361898 364226
rect 361718 364046 361774 364102
rect 361842 364046 361898 364102
rect 361718 363922 361774 363978
rect 361842 363922 361898 363978
rect 392438 364294 392494 364350
rect 392562 364294 392618 364350
rect 392438 364170 392494 364226
rect 392562 364170 392618 364226
rect 392438 364046 392494 364102
rect 392562 364046 392618 364102
rect 392438 363922 392494 363978
rect 392562 363922 392618 363978
rect 423158 364294 423214 364350
rect 423282 364294 423338 364350
rect 423158 364170 423214 364226
rect 423282 364170 423338 364226
rect 423158 364046 423214 364102
rect 423282 364046 423338 364102
rect 423158 363922 423214 363978
rect 423282 363922 423338 363978
rect 453878 364294 453934 364350
rect 454002 364294 454058 364350
rect 453878 364170 453934 364226
rect 454002 364170 454058 364226
rect 453878 364046 453934 364102
rect 454002 364046 454058 364102
rect 453878 363922 453934 363978
rect 454002 363922 454058 363978
rect 484598 364294 484654 364350
rect 484722 364294 484778 364350
rect 484598 364170 484654 364226
rect 484722 364170 484778 364226
rect 484598 364046 484654 364102
rect 484722 364046 484778 364102
rect 484598 363922 484654 363978
rect 484722 363922 484778 363978
rect 515318 364294 515374 364350
rect 515442 364294 515498 364350
rect 515318 364170 515374 364226
rect 515442 364170 515498 364226
rect 515318 364046 515374 364102
rect 515442 364046 515498 364102
rect 515318 363922 515374 363978
rect 515442 363922 515498 363978
rect 546038 364294 546094 364350
rect 546162 364294 546218 364350
rect 546038 364170 546094 364226
rect 546162 364170 546218 364226
rect 546038 364046 546094 364102
rect 546162 364046 546218 364102
rect 546038 363922 546094 363978
rect 546162 363922 546218 363978
rect 561250 364294 561306 364350
rect 561374 364294 561430 364350
rect 561498 364294 561554 364350
rect 561622 364294 561678 364350
rect 561250 364170 561306 364226
rect 561374 364170 561430 364226
rect 561498 364170 561554 364226
rect 561622 364170 561678 364226
rect 561250 364046 561306 364102
rect 561374 364046 561430 364102
rect 561498 364046 561554 364102
rect 561622 364046 561678 364102
rect 561250 363922 561306 363978
rect 561374 363922 561430 363978
rect 561498 363922 561554 363978
rect 561622 363922 561678 363978
rect 131318 352294 131374 352350
rect 131442 352294 131498 352350
rect 131318 352170 131374 352226
rect 131442 352170 131498 352226
rect 131318 352046 131374 352102
rect 131442 352046 131498 352102
rect 131318 351922 131374 351978
rect 131442 351922 131498 351978
rect 162038 352294 162094 352350
rect 162162 352294 162218 352350
rect 162038 352170 162094 352226
rect 162162 352170 162218 352226
rect 162038 352046 162094 352102
rect 162162 352046 162218 352102
rect 162038 351922 162094 351978
rect 162162 351922 162218 351978
rect 192758 352294 192814 352350
rect 192882 352294 192938 352350
rect 192758 352170 192814 352226
rect 192882 352170 192938 352226
rect 192758 352046 192814 352102
rect 192882 352046 192938 352102
rect 192758 351922 192814 351978
rect 192882 351922 192938 351978
rect 223478 352294 223534 352350
rect 223602 352294 223658 352350
rect 223478 352170 223534 352226
rect 223602 352170 223658 352226
rect 223478 352046 223534 352102
rect 223602 352046 223658 352102
rect 223478 351922 223534 351978
rect 223602 351922 223658 351978
rect 254198 352294 254254 352350
rect 254322 352294 254378 352350
rect 254198 352170 254254 352226
rect 254322 352170 254378 352226
rect 254198 352046 254254 352102
rect 254322 352046 254378 352102
rect 254198 351922 254254 351978
rect 254322 351922 254378 351978
rect 284918 352294 284974 352350
rect 285042 352294 285098 352350
rect 284918 352170 284974 352226
rect 285042 352170 285098 352226
rect 284918 352046 284974 352102
rect 285042 352046 285098 352102
rect 284918 351922 284974 351978
rect 285042 351922 285098 351978
rect 315638 352294 315694 352350
rect 315762 352294 315818 352350
rect 315638 352170 315694 352226
rect 315762 352170 315818 352226
rect 315638 352046 315694 352102
rect 315762 352046 315818 352102
rect 315638 351922 315694 351978
rect 315762 351922 315818 351978
rect 346358 352294 346414 352350
rect 346482 352294 346538 352350
rect 346358 352170 346414 352226
rect 346482 352170 346538 352226
rect 346358 352046 346414 352102
rect 346482 352046 346538 352102
rect 346358 351922 346414 351978
rect 346482 351922 346538 351978
rect 377078 352294 377134 352350
rect 377202 352294 377258 352350
rect 377078 352170 377134 352226
rect 377202 352170 377258 352226
rect 377078 352046 377134 352102
rect 377202 352046 377258 352102
rect 377078 351922 377134 351978
rect 377202 351922 377258 351978
rect 407798 352294 407854 352350
rect 407922 352294 407978 352350
rect 407798 352170 407854 352226
rect 407922 352170 407978 352226
rect 407798 352046 407854 352102
rect 407922 352046 407978 352102
rect 407798 351922 407854 351978
rect 407922 351922 407978 351978
rect 438518 352294 438574 352350
rect 438642 352294 438698 352350
rect 438518 352170 438574 352226
rect 438642 352170 438698 352226
rect 438518 352046 438574 352102
rect 438642 352046 438698 352102
rect 438518 351922 438574 351978
rect 438642 351922 438698 351978
rect 469238 352294 469294 352350
rect 469362 352294 469418 352350
rect 469238 352170 469294 352226
rect 469362 352170 469418 352226
rect 469238 352046 469294 352102
rect 469362 352046 469418 352102
rect 469238 351922 469294 351978
rect 469362 351922 469418 351978
rect 499958 352294 500014 352350
rect 500082 352294 500138 352350
rect 499958 352170 500014 352226
rect 500082 352170 500138 352226
rect 499958 352046 500014 352102
rect 500082 352046 500138 352102
rect 499958 351922 500014 351978
rect 500082 351922 500138 351978
rect 530678 352294 530734 352350
rect 530802 352294 530858 352350
rect 530678 352170 530734 352226
rect 530802 352170 530858 352226
rect 530678 352046 530734 352102
rect 530802 352046 530858 352102
rect 530678 351922 530734 351978
rect 530802 351922 530858 351978
rect 111250 346294 111306 346350
rect 111374 346294 111430 346350
rect 111498 346294 111554 346350
rect 111622 346294 111678 346350
rect 111250 346170 111306 346226
rect 111374 346170 111430 346226
rect 111498 346170 111554 346226
rect 111622 346170 111678 346226
rect 111250 346046 111306 346102
rect 111374 346046 111430 346102
rect 111498 346046 111554 346102
rect 111622 346046 111678 346102
rect 111250 345922 111306 345978
rect 111374 345922 111430 345978
rect 111498 345922 111554 345978
rect 111622 345922 111678 345978
rect 96970 334294 97026 334350
rect 97094 334294 97150 334350
rect 97218 334294 97274 334350
rect 97342 334294 97398 334350
rect 96970 334170 97026 334226
rect 97094 334170 97150 334226
rect 97218 334170 97274 334226
rect 97342 334170 97398 334226
rect 96970 334046 97026 334102
rect 97094 334046 97150 334102
rect 97218 334046 97274 334102
rect 97342 334046 97398 334102
rect 96970 333922 97026 333978
rect 97094 333922 97150 333978
rect 97218 333922 97274 333978
rect 97342 333922 97398 333978
rect 100598 334294 100654 334350
rect 100722 334294 100778 334350
rect 100598 334170 100654 334226
rect 100722 334170 100778 334226
rect 100598 334046 100654 334102
rect 100722 334046 100778 334102
rect 100598 333922 100654 333978
rect 100722 333922 100778 333978
rect 115958 346294 116014 346350
rect 116082 346294 116138 346350
rect 115958 346170 116014 346226
rect 116082 346170 116138 346226
rect 115958 346046 116014 346102
rect 116082 346046 116138 346102
rect 115958 345922 116014 345978
rect 116082 345922 116138 345978
rect 146678 346294 146734 346350
rect 146802 346294 146858 346350
rect 146678 346170 146734 346226
rect 146802 346170 146858 346226
rect 146678 346046 146734 346102
rect 146802 346046 146858 346102
rect 146678 345922 146734 345978
rect 146802 345922 146858 345978
rect 177398 346294 177454 346350
rect 177522 346294 177578 346350
rect 177398 346170 177454 346226
rect 177522 346170 177578 346226
rect 177398 346046 177454 346102
rect 177522 346046 177578 346102
rect 177398 345922 177454 345978
rect 177522 345922 177578 345978
rect 208118 346294 208174 346350
rect 208242 346294 208298 346350
rect 208118 346170 208174 346226
rect 208242 346170 208298 346226
rect 208118 346046 208174 346102
rect 208242 346046 208298 346102
rect 208118 345922 208174 345978
rect 208242 345922 208298 345978
rect 238838 346294 238894 346350
rect 238962 346294 239018 346350
rect 238838 346170 238894 346226
rect 238962 346170 239018 346226
rect 238838 346046 238894 346102
rect 238962 346046 239018 346102
rect 238838 345922 238894 345978
rect 238962 345922 239018 345978
rect 269558 346294 269614 346350
rect 269682 346294 269738 346350
rect 269558 346170 269614 346226
rect 269682 346170 269738 346226
rect 269558 346046 269614 346102
rect 269682 346046 269738 346102
rect 269558 345922 269614 345978
rect 269682 345922 269738 345978
rect 300278 346294 300334 346350
rect 300402 346294 300458 346350
rect 300278 346170 300334 346226
rect 300402 346170 300458 346226
rect 300278 346046 300334 346102
rect 300402 346046 300458 346102
rect 300278 345922 300334 345978
rect 300402 345922 300458 345978
rect 330998 346294 331054 346350
rect 331122 346294 331178 346350
rect 330998 346170 331054 346226
rect 331122 346170 331178 346226
rect 330998 346046 331054 346102
rect 331122 346046 331178 346102
rect 330998 345922 331054 345978
rect 331122 345922 331178 345978
rect 361718 346294 361774 346350
rect 361842 346294 361898 346350
rect 361718 346170 361774 346226
rect 361842 346170 361898 346226
rect 361718 346046 361774 346102
rect 361842 346046 361898 346102
rect 361718 345922 361774 345978
rect 361842 345922 361898 345978
rect 392438 346294 392494 346350
rect 392562 346294 392618 346350
rect 392438 346170 392494 346226
rect 392562 346170 392618 346226
rect 392438 346046 392494 346102
rect 392562 346046 392618 346102
rect 392438 345922 392494 345978
rect 392562 345922 392618 345978
rect 423158 346294 423214 346350
rect 423282 346294 423338 346350
rect 423158 346170 423214 346226
rect 423282 346170 423338 346226
rect 423158 346046 423214 346102
rect 423282 346046 423338 346102
rect 423158 345922 423214 345978
rect 423282 345922 423338 345978
rect 453878 346294 453934 346350
rect 454002 346294 454058 346350
rect 453878 346170 453934 346226
rect 454002 346170 454058 346226
rect 453878 346046 453934 346102
rect 454002 346046 454058 346102
rect 453878 345922 453934 345978
rect 454002 345922 454058 345978
rect 484598 346294 484654 346350
rect 484722 346294 484778 346350
rect 484598 346170 484654 346226
rect 484722 346170 484778 346226
rect 484598 346046 484654 346102
rect 484722 346046 484778 346102
rect 484598 345922 484654 345978
rect 484722 345922 484778 345978
rect 515318 346294 515374 346350
rect 515442 346294 515498 346350
rect 515318 346170 515374 346226
rect 515442 346170 515498 346226
rect 515318 346046 515374 346102
rect 515442 346046 515498 346102
rect 515318 345922 515374 345978
rect 515442 345922 515498 345978
rect 546038 346294 546094 346350
rect 546162 346294 546218 346350
rect 546038 346170 546094 346226
rect 546162 346170 546218 346226
rect 546038 346046 546094 346102
rect 546162 346046 546218 346102
rect 546038 345922 546094 345978
rect 546162 345922 546218 345978
rect 561250 346294 561306 346350
rect 561374 346294 561430 346350
rect 561498 346294 561554 346350
rect 561622 346294 561678 346350
rect 561250 346170 561306 346226
rect 561374 346170 561430 346226
rect 561498 346170 561554 346226
rect 561622 346170 561678 346226
rect 561250 346046 561306 346102
rect 561374 346046 561430 346102
rect 561498 346046 561554 346102
rect 561622 346046 561678 346102
rect 561250 345922 561306 345978
rect 561374 345922 561430 345978
rect 561498 345922 561554 345978
rect 561622 345922 561678 345978
rect 131318 334294 131374 334350
rect 131442 334294 131498 334350
rect 131318 334170 131374 334226
rect 131442 334170 131498 334226
rect 131318 334046 131374 334102
rect 131442 334046 131498 334102
rect 131318 333922 131374 333978
rect 131442 333922 131498 333978
rect 162038 334294 162094 334350
rect 162162 334294 162218 334350
rect 162038 334170 162094 334226
rect 162162 334170 162218 334226
rect 162038 334046 162094 334102
rect 162162 334046 162218 334102
rect 162038 333922 162094 333978
rect 162162 333922 162218 333978
rect 192758 334294 192814 334350
rect 192882 334294 192938 334350
rect 192758 334170 192814 334226
rect 192882 334170 192938 334226
rect 192758 334046 192814 334102
rect 192882 334046 192938 334102
rect 192758 333922 192814 333978
rect 192882 333922 192938 333978
rect 223478 334294 223534 334350
rect 223602 334294 223658 334350
rect 223478 334170 223534 334226
rect 223602 334170 223658 334226
rect 223478 334046 223534 334102
rect 223602 334046 223658 334102
rect 223478 333922 223534 333978
rect 223602 333922 223658 333978
rect 254198 334294 254254 334350
rect 254322 334294 254378 334350
rect 254198 334170 254254 334226
rect 254322 334170 254378 334226
rect 254198 334046 254254 334102
rect 254322 334046 254378 334102
rect 254198 333922 254254 333978
rect 254322 333922 254378 333978
rect 284918 334294 284974 334350
rect 285042 334294 285098 334350
rect 284918 334170 284974 334226
rect 285042 334170 285098 334226
rect 284918 334046 284974 334102
rect 285042 334046 285098 334102
rect 284918 333922 284974 333978
rect 285042 333922 285098 333978
rect 315638 334294 315694 334350
rect 315762 334294 315818 334350
rect 315638 334170 315694 334226
rect 315762 334170 315818 334226
rect 315638 334046 315694 334102
rect 315762 334046 315818 334102
rect 315638 333922 315694 333978
rect 315762 333922 315818 333978
rect 346358 334294 346414 334350
rect 346482 334294 346538 334350
rect 346358 334170 346414 334226
rect 346482 334170 346538 334226
rect 346358 334046 346414 334102
rect 346482 334046 346538 334102
rect 346358 333922 346414 333978
rect 346482 333922 346538 333978
rect 377078 334294 377134 334350
rect 377202 334294 377258 334350
rect 377078 334170 377134 334226
rect 377202 334170 377258 334226
rect 377078 334046 377134 334102
rect 377202 334046 377258 334102
rect 377078 333922 377134 333978
rect 377202 333922 377258 333978
rect 407798 334294 407854 334350
rect 407922 334294 407978 334350
rect 407798 334170 407854 334226
rect 407922 334170 407978 334226
rect 407798 334046 407854 334102
rect 407922 334046 407978 334102
rect 407798 333922 407854 333978
rect 407922 333922 407978 333978
rect 438518 334294 438574 334350
rect 438642 334294 438698 334350
rect 438518 334170 438574 334226
rect 438642 334170 438698 334226
rect 438518 334046 438574 334102
rect 438642 334046 438698 334102
rect 438518 333922 438574 333978
rect 438642 333922 438698 333978
rect 469238 334294 469294 334350
rect 469362 334294 469418 334350
rect 469238 334170 469294 334226
rect 469362 334170 469418 334226
rect 469238 334046 469294 334102
rect 469362 334046 469418 334102
rect 469238 333922 469294 333978
rect 469362 333922 469418 333978
rect 499958 334294 500014 334350
rect 500082 334294 500138 334350
rect 499958 334170 500014 334226
rect 500082 334170 500138 334226
rect 499958 334046 500014 334102
rect 500082 334046 500138 334102
rect 499958 333922 500014 333978
rect 500082 333922 500138 333978
rect 530678 334294 530734 334350
rect 530802 334294 530858 334350
rect 530678 334170 530734 334226
rect 530802 334170 530858 334226
rect 530678 334046 530734 334102
rect 530802 334046 530858 334102
rect 530678 333922 530734 333978
rect 530802 333922 530858 333978
rect 111250 328294 111306 328350
rect 111374 328294 111430 328350
rect 111498 328294 111554 328350
rect 111622 328294 111678 328350
rect 111250 328170 111306 328226
rect 111374 328170 111430 328226
rect 111498 328170 111554 328226
rect 111622 328170 111678 328226
rect 111250 328046 111306 328102
rect 111374 328046 111430 328102
rect 111498 328046 111554 328102
rect 111622 328046 111678 328102
rect 111250 327922 111306 327978
rect 111374 327922 111430 327978
rect 111498 327922 111554 327978
rect 111622 327922 111678 327978
rect 96970 316294 97026 316350
rect 97094 316294 97150 316350
rect 97218 316294 97274 316350
rect 97342 316294 97398 316350
rect 96970 316170 97026 316226
rect 97094 316170 97150 316226
rect 97218 316170 97274 316226
rect 97342 316170 97398 316226
rect 96970 316046 97026 316102
rect 97094 316046 97150 316102
rect 97218 316046 97274 316102
rect 97342 316046 97398 316102
rect 96970 315922 97026 315978
rect 97094 315922 97150 315978
rect 97218 315922 97274 315978
rect 97342 315922 97398 315978
rect 100598 316294 100654 316350
rect 100722 316294 100778 316350
rect 100598 316170 100654 316226
rect 100722 316170 100778 316226
rect 100598 316046 100654 316102
rect 100722 316046 100778 316102
rect 100598 315922 100654 315978
rect 100722 315922 100778 315978
rect 115958 328294 116014 328350
rect 116082 328294 116138 328350
rect 115958 328170 116014 328226
rect 116082 328170 116138 328226
rect 115958 328046 116014 328102
rect 116082 328046 116138 328102
rect 115958 327922 116014 327978
rect 116082 327922 116138 327978
rect 146678 328294 146734 328350
rect 146802 328294 146858 328350
rect 146678 328170 146734 328226
rect 146802 328170 146858 328226
rect 146678 328046 146734 328102
rect 146802 328046 146858 328102
rect 146678 327922 146734 327978
rect 146802 327922 146858 327978
rect 177398 328294 177454 328350
rect 177522 328294 177578 328350
rect 177398 328170 177454 328226
rect 177522 328170 177578 328226
rect 177398 328046 177454 328102
rect 177522 328046 177578 328102
rect 177398 327922 177454 327978
rect 177522 327922 177578 327978
rect 208118 328294 208174 328350
rect 208242 328294 208298 328350
rect 208118 328170 208174 328226
rect 208242 328170 208298 328226
rect 208118 328046 208174 328102
rect 208242 328046 208298 328102
rect 208118 327922 208174 327978
rect 208242 327922 208298 327978
rect 238838 328294 238894 328350
rect 238962 328294 239018 328350
rect 238838 328170 238894 328226
rect 238962 328170 239018 328226
rect 238838 328046 238894 328102
rect 238962 328046 239018 328102
rect 238838 327922 238894 327978
rect 238962 327922 239018 327978
rect 269558 328294 269614 328350
rect 269682 328294 269738 328350
rect 269558 328170 269614 328226
rect 269682 328170 269738 328226
rect 269558 328046 269614 328102
rect 269682 328046 269738 328102
rect 269558 327922 269614 327978
rect 269682 327922 269738 327978
rect 300278 328294 300334 328350
rect 300402 328294 300458 328350
rect 300278 328170 300334 328226
rect 300402 328170 300458 328226
rect 300278 328046 300334 328102
rect 300402 328046 300458 328102
rect 300278 327922 300334 327978
rect 300402 327922 300458 327978
rect 330998 328294 331054 328350
rect 331122 328294 331178 328350
rect 330998 328170 331054 328226
rect 331122 328170 331178 328226
rect 330998 328046 331054 328102
rect 331122 328046 331178 328102
rect 330998 327922 331054 327978
rect 331122 327922 331178 327978
rect 361718 328294 361774 328350
rect 361842 328294 361898 328350
rect 361718 328170 361774 328226
rect 361842 328170 361898 328226
rect 361718 328046 361774 328102
rect 361842 328046 361898 328102
rect 361718 327922 361774 327978
rect 361842 327922 361898 327978
rect 392438 328294 392494 328350
rect 392562 328294 392618 328350
rect 392438 328170 392494 328226
rect 392562 328170 392618 328226
rect 392438 328046 392494 328102
rect 392562 328046 392618 328102
rect 392438 327922 392494 327978
rect 392562 327922 392618 327978
rect 423158 328294 423214 328350
rect 423282 328294 423338 328350
rect 423158 328170 423214 328226
rect 423282 328170 423338 328226
rect 423158 328046 423214 328102
rect 423282 328046 423338 328102
rect 423158 327922 423214 327978
rect 423282 327922 423338 327978
rect 453878 328294 453934 328350
rect 454002 328294 454058 328350
rect 453878 328170 453934 328226
rect 454002 328170 454058 328226
rect 453878 328046 453934 328102
rect 454002 328046 454058 328102
rect 453878 327922 453934 327978
rect 454002 327922 454058 327978
rect 484598 328294 484654 328350
rect 484722 328294 484778 328350
rect 484598 328170 484654 328226
rect 484722 328170 484778 328226
rect 484598 328046 484654 328102
rect 484722 328046 484778 328102
rect 484598 327922 484654 327978
rect 484722 327922 484778 327978
rect 515318 328294 515374 328350
rect 515442 328294 515498 328350
rect 515318 328170 515374 328226
rect 515442 328170 515498 328226
rect 515318 328046 515374 328102
rect 515442 328046 515498 328102
rect 515318 327922 515374 327978
rect 515442 327922 515498 327978
rect 546038 328294 546094 328350
rect 546162 328294 546218 328350
rect 546038 328170 546094 328226
rect 546162 328170 546218 328226
rect 546038 328046 546094 328102
rect 546162 328046 546218 328102
rect 546038 327922 546094 327978
rect 546162 327922 546218 327978
rect 561250 328294 561306 328350
rect 561374 328294 561430 328350
rect 561498 328294 561554 328350
rect 561622 328294 561678 328350
rect 561250 328170 561306 328226
rect 561374 328170 561430 328226
rect 561498 328170 561554 328226
rect 561622 328170 561678 328226
rect 561250 328046 561306 328102
rect 561374 328046 561430 328102
rect 561498 328046 561554 328102
rect 561622 328046 561678 328102
rect 561250 327922 561306 327978
rect 561374 327922 561430 327978
rect 561498 327922 561554 327978
rect 561622 327922 561678 327978
rect 131318 316294 131374 316350
rect 131442 316294 131498 316350
rect 131318 316170 131374 316226
rect 131442 316170 131498 316226
rect 131318 316046 131374 316102
rect 131442 316046 131498 316102
rect 131318 315922 131374 315978
rect 131442 315922 131498 315978
rect 162038 316294 162094 316350
rect 162162 316294 162218 316350
rect 162038 316170 162094 316226
rect 162162 316170 162218 316226
rect 162038 316046 162094 316102
rect 162162 316046 162218 316102
rect 162038 315922 162094 315978
rect 162162 315922 162218 315978
rect 192758 316294 192814 316350
rect 192882 316294 192938 316350
rect 192758 316170 192814 316226
rect 192882 316170 192938 316226
rect 192758 316046 192814 316102
rect 192882 316046 192938 316102
rect 192758 315922 192814 315978
rect 192882 315922 192938 315978
rect 223478 316294 223534 316350
rect 223602 316294 223658 316350
rect 223478 316170 223534 316226
rect 223602 316170 223658 316226
rect 223478 316046 223534 316102
rect 223602 316046 223658 316102
rect 223478 315922 223534 315978
rect 223602 315922 223658 315978
rect 254198 316294 254254 316350
rect 254322 316294 254378 316350
rect 254198 316170 254254 316226
rect 254322 316170 254378 316226
rect 254198 316046 254254 316102
rect 254322 316046 254378 316102
rect 254198 315922 254254 315978
rect 254322 315922 254378 315978
rect 284918 316294 284974 316350
rect 285042 316294 285098 316350
rect 284918 316170 284974 316226
rect 285042 316170 285098 316226
rect 284918 316046 284974 316102
rect 285042 316046 285098 316102
rect 284918 315922 284974 315978
rect 285042 315922 285098 315978
rect 315638 316294 315694 316350
rect 315762 316294 315818 316350
rect 315638 316170 315694 316226
rect 315762 316170 315818 316226
rect 315638 316046 315694 316102
rect 315762 316046 315818 316102
rect 315638 315922 315694 315978
rect 315762 315922 315818 315978
rect 346358 316294 346414 316350
rect 346482 316294 346538 316350
rect 346358 316170 346414 316226
rect 346482 316170 346538 316226
rect 346358 316046 346414 316102
rect 346482 316046 346538 316102
rect 346358 315922 346414 315978
rect 346482 315922 346538 315978
rect 377078 316294 377134 316350
rect 377202 316294 377258 316350
rect 377078 316170 377134 316226
rect 377202 316170 377258 316226
rect 377078 316046 377134 316102
rect 377202 316046 377258 316102
rect 377078 315922 377134 315978
rect 377202 315922 377258 315978
rect 407798 316294 407854 316350
rect 407922 316294 407978 316350
rect 407798 316170 407854 316226
rect 407922 316170 407978 316226
rect 407798 316046 407854 316102
rect 407922 316046 407978 316102
rect 407798 315922 407854 315978
rect 407922 315922 407978 315978
rect 438518 316294 438574 316350
rect 438642 316294 438698 316350
rect 438518 316170 438574 316226
rect 438642 316170 438698 316226
rect 438518 316046 438574 316102
rect 438642 316046 438698 316102
rect 438518 315922 438574 315978
rect 438642 315922 438698 315978
rect 469238 316294 469294 316350
rect 469362 316294 469418 316350
rect 469238 316170 469294 316226
rect 469362 316170 469418 316226
rect 469238 316046 469294 316102
rect 469362 316046 469418 316102
rect 469238 315922 469294 315978
rect 469362 315922 469418 315978
rect 499958 316294 500014 316350
rect 500082 316294 500138 316350
rect 499958 316170 500014 316226
rect 500082 316170 500138 316226
rect 499958 316046 500014 316102
rect 500082 316046 500138 316102
rect 499958 315922 500014 315978
rect 500082 315922 500138 315978
rect 530678 316294 530734 316350
rect 530802 316294 530858 316350
rect 530678 316170 530734 316226
rect 530802 316170 530858 316226
rect 530678 316046 530734 316102
rect 530802 316046 530858 316102
rect 530678 315922 530734 315978
rect 530802 315922 530858 315978
rect 111250 310294 111306 310350
rect 111374 310294 111430 310350
rect 111498 310294 111554 310350
rect 111622 310294 111678 310350
rect 111250 310170 111306 310226
rect 111374 310170 111430 310226
rect 111498 310170 111554 310226
rect 111622 310170 111678 310226
rect 111250 310046 111306 310102
rect 111374 310046 111430 310102
rect 111498 310046 111554 310102
rect 111622 310046 111678 310102
rect 111250 309922 111306 309978
rect 111374 309922 111430 309978
rect 111498 309922 111554 309978
rect 111622 309922 111678 309978
rect 96970 298294 97026 298350
rect 97094 298294 97150 298350
rect 97218 298294 97274 298350
rect 97342 298294 97398 298350
rect 96970 298170 97026 298226
rect 97094 298170 97150 298226
rect 97218 298170 97274 298226
rect 97342 298170 97398 298226
rect 96970 298046 97026 298102
rect 97094 298046 97150 298102
rect 97218 298046 97274 298102
rect 97342 298046 97398 298102
rect 96970 297922 97026 297978
rect 97094 297922 97150 297978
rect 97218 297922 97274 297978
rect 97342 297922 97398 297978
rect 100598 298294 100654 298350
rect 100722 298294 100778 298350
rect 100598 298170 100654 298226
rect 100722 298170 100778 298226
rect 100598 298046 100654 298102
rect 100722 298046 100778 298102
rect 100598 297922 100654 297978
rect 100722 297922 100778 297978
rect 115958 310294 116014 310350
rect 116082 310294 116138 310350
rect 115958 310170 116014 310226
rect 116082 310170 116138 310226
rect 115958 310046 116014 310102
rect 116082 310046 116138 310102
rect 115958 309922 116014 309978
rect 116082 309922 116138 309978
rect 146678 310294 146734 310350
rect 146802 310294 146858 310350
rect 146678 310170 146734 310226
rect 146802 310170 146858 310226
rect 146678 310046 146734 310102
rect 146802 310046 146858 310102
rect 146678 309922 146734 309978
rect 146802 309922 146858 309978
rect 177398 310294 177454 310350
rect 177522 310294 177578 310350
rect 177398 310170 177454 310226
rect 177522 310170 177578 310226
rect 177398 310046 177454 310102
rect 177522 310046 177578 310102
rect 177398 309922 177454 309978
rect 177522 309922 177578 309978
rect 208118 310294 208174 310350
rect 208242 310294 208298 310350
rect 208118 310170 208174 310226
rect 208242 310170 208298 310226
rect 208118 310046 208174 310102
rect 208242 310046 208298 310102
rect 208118 309922 208174 309978
rect 208242 309922 208298 309978
rect 238838 310294 238894 310350
rect 238962 310294 239018 310350
rect 238838 310170 238894 310226
rect 238962 310170 239018 310226
rect 238838 310046 238894 310102
rect 238962 310046 239018 310102
rect 238838 309922 238894 309978
rect 238962 309922 239018 309978
rect 269558 310294 269614 310350
rect 269682 310294 269738 310350
rect 269558 310170 269614 310226
rect 269682 310170 269738 310226
rect 269558 310046 269614 310102
rect 269682 310046 269738 310102
rect 269558 309922 269614 309978
rect 269682 309922 269738 309978
rect 300278 310294 300334 310350
rect 300402 310294 300458 310350
rect 300278 310170 300334 310226
rect 300402 310170 300458 310226
rect 300278 310046 300334 310102
rect 300402 310046 300458 310102
rect 300278 309922 300334 309978
rect 300402 309922 300458 309978
rect 330998 310294 331054 310350
rect 331122 310294 331178 310350
rect 330998 310170 331054 310226
rect 331122 310170 331178 310226
rect 330998 310046 331054 310102
rect 331122 310046 331178 310102
rect 330998 309922 331054 309978
rect 331122 309922 331178 309978
rect 361718 310294 361774 310350
rect 361842 310294 361898 310350
rect 361718 310170 361774 310226
rect 361842 310170 361898 310226
rect 361718 310046 361774 310102
rect 361842 310046 361898 310102
rect 361718 309922 361774 309978
rect 361842 309922 361898 309978
rect 392438 310294 392494 310350
rect 392562 310294 392618 310350
rect 392438 310170 392494 310226
rect 392562 310170 392618 310226
rect 392438 310046 392494 310102
rect 392562 310046 392618 310102
rect 392438 309922 392494 309978
rect 392562 309922 392618 309978
rect 423158 310294 423214 310350
rect 423282 310294 423338 310350
rect 423158 310170 423214 310226
rect 423282 310170 423338 310226
rect 423158 310046 423214 310102
rect 423282 310046 423338 310102
rect 423158 309922 423214 309978
rect 423282 309922 423338 309978
rect 453878 310294 453934 310350
rect 454002 310294 454058 310350
rect 453878 310170 453934 310226
rect 454002 310170 454058 310226
rect 453878 310046 453934 310102
rect 454002 310046 454058 310102
rect 453878 309922 453934 309978
rect 454002 309922 454058 309978
rect 484598 310294 484654 310350
rect 484722 310294 484778 310350
rect 484598 310170 484654 310226
rect 484722 310170 484778 310226
rect 484598 310046 484654 310102
rect 484722 310046 484778 310102
rect 484598 309922 484654 309978
rect 484722 309922 484778 309978
rect 515318 310294 515374 310350
rect 515442 310294 515498 310350
rect 515318 310170 515374 310226
rect 515442 310170 515498 310226
rect 515318 310046 515374 310102
rect 515442 310046 515498 310102
rect 515318 309922 515374 309978
rect 515442 309922 515498 309978
rect 546038 310294 546094 310350
rect 546162 310294 546218 310350
rect 546038 310170 546094 310226
rect 546162 310170 546218 310226
rect 546038 310046 546094 310102
rect 546162 310046 546218 310102
rect 546038 309922 546094 309978
rect 546162 309922 546218 309978
rect 561250 310294 561306 310350
rect 561374 310294 561430 310350
rect 561498 310294 561554 310350
rect 561622 310294 561678 310350
rect 561250 310170 561306 310226
rect 561374 310170 561430 310226
rect 561498 310170 561554 310226
rect 561622 310170 561678 310226
rect 561250 310046 561306 310102
rect 561374 310046 561430 310102
rect 561498 310046 561554 310102
rect 561622 310046 561678 310102
rect 561250 309922 561306 309978
rect 561374 309922 561430 309978
rect 561498 309922 561554 309978
rect 561622 309922 561678 309978
rect 131318 298294 131374 298350
rect 131442 298294 131498 298350
rect 131318 298170 131374 298226
rect 131442 298170 131498 298226
rect 131318 298046 131374 298102
rect 131442 298046 131498 298102
rect 131318 297922 131374 297978
rect 131442 297922 131498 297978
rect 162038 298294 162094 298350
rect 162162 298294 162218 298350
rect 162038 298170 162094 298226
rect 162162 298170 162218 298226
rect 162038 298046 162094 298102
rect 162162 298046 162218 298102
rect 162038 297922 162094 297978
rect 162162 297922 162218 297978
rect 192758 298294 192814 298350
rect 192882 298294 192938 298350
rect 192758 298170 192814 298226
rect 192882 298170 192938 298226
rect 192758 298046 192814 298102
rect 192882 298046 192938 298102
rect 192758 297922 192814 297978
rect 192882 297922 192938 297978
rect 223478 298294 223534 298350
rect 223602 298294 223658 298350
rect 223478 298170 223534 298226
rect 223602 298170 223658 298226
rect 223478 298046 223534 298102
rect 223602 298046 223658 298102
rect 223478 297922 223534 297978
rect 223602 297922 223658 297978
rect 254198 298294 254254 298350
rect 254322 298294 254378 298350
rect 254198 298170 254254 298226
rect 254322 298170 254378 298226
rect 254198 298046 254254 298102
rect 254322 298046 254378 298102
rect 254198 297922 254254 297978
rect 254322 297922 254378 297978
rect 284918 298294 284974 298350
rect 285042 298294 285098 298350
rect 284918 298170 284974 298226
rect 285042 298170 285098 298226
rect 284918 298046 284974 298102
rect 285042 298046 285098 298102
rect 284918 297922 284974 297978
rect 285042 297922 285098 297978
rect 315638 298294 315694 298350
rect 315762 298294 315818 298350
rect 315638 298170 315694 298226
rect 315762 298170 315818 298226
rect 315638 298046 315694 298102
rect 315762 298046 315818 298102
rect 315638 297922 315694 297978
rect 315762 297922 315818 297978
rect 346358 298294 346414 298350
rect 346482 298294 346538 298350
rect 346358 298170 346414 298226
rect 346482 298170 346538 298226
rect 346358 298046 346414 298102
rect 346482 298046 346538 298102
rect 346358 297922 346414 297978
rect 346482 297922 346538 297978
rect 377078 298294 377134 298350
rect 377202 298294 377258 298350
rect 377078 298170 377134 298226
rect 377202 298170 377258 298226
rect 377078 298046 377134 298102
rect 377202 298046 377258 298102
rect 377078 297922 377134 297978
rect 377202 297922 377258 297978
rect 407798 298294 407854 298350
rect 407922 298294 407978 298350
rect 407798 298170 407854 298226
rect 407922 298170 407978 298226
rect 407798 298046 407854 298102
rect 407922 298046 407978 298102
rect 407798 297922 407854 297978
rect 407922 297922 407978 297978
rect 438518 298294 438574 298350
rect 438642 298294 438698 298350
rect 438518 298170 438574 298226
rect 438642 298170 438698 298226
rect 438518 298046 438574 298102
rect 438642 298046 438698 298102
rect 438518 297922 438574 297978
rect 438642 297922 438698 297978
rect 469238 298294 469294 298350
rect 469362 298294 469418 298350
rect 469238 298170 469294 298226
rect 469362 298170 469418 298226
rect 469238 298046 469294 298102
rect 469362 298046 469418 298102
rect 469238 297922 469294 297978
rect 469362 297922 469418 297978
rect 499958 298294 500014 298350
rect 500082 298294 500138 298350
rect 499958 298170 500014 298226
rect 500082 298170 500138 298226
rect 499958 298046 500014 298102
rect 500082 298046 500138 298102
rect 499958 297922 500014 297978
rect 500082 297922 500138 297978
rect 530678 298294 530734 298350
rect 530802 298294 530858 298350
rect 530678 298170 530734 298226
rect 530802 298170 530858 298226
rect 530678 298046 530734 298102
rect 530802 298046 530858 298102
rect 530678 297922 530734 297978
rect 530802 297922 530858 297978
rect 111250 292294 111306 292350
rect 111374 292294 111430 292350
rect 111498 292294 111554 292350
rect 111622 292294 111678 292350
rect 111250 292170 111306 292226
rect 111374 292170 111430 292226
rect 111498 292170 111554 292226
rect 111622 292170 111678 292226
rect 111250 292046 111306 292102
rect 111374 292046 111430 292102
rect 111498 292046 111554 292102
rect 111622 292046 111678 292102
rect 111250 291922 111306 291978
rect 111374 291922 111430 291978
rect 111498 291922 111554 291978
rect 111622 291922 111678 291978
rect 96970 280294 97026 280350
rect 97094 280294 97150 280350
rect 97218 280294 97274 280350
rect 97342 280294 97398 280350
rect 96970 280170 97026 280226
rect 97094 280170 97150 280226
rect 97218 280170 97274 280226
rect 97342 280170 97398 280226
rect 96970 280046 97026 280102
rect 97094 280046 97150 280102
rect 97218 280046 97274 280102
rect 97342 280046 97398 280102
rect 96970 279922 97026 279978
rect 97094 279922 97150 279978
rect 97218 279922 97274 279978
rect 97342 279922 97398 279978
rect 100598 280294 100654 280350
rect 100722 280294 100778 280350
rect 100598 280170 100654 280226
rect 100722 280170 100778 280226
rect 100598 280046 100654 280102
rect 100722 280046 100778 280102
rect 100598 279922 100654 279978
rect 100722 279922 100778 279978
rect 115958 292294 116014 292350
rect 116082 292294 116138 292350
rect 115958 292170 116014 292226
rect 116082 292170 116138 292226
rect 115958 292046 116014 292102
rect 116082 292046 116138 292102
rect 115958 291922 116014 291978
rect 116082 291922 116138 291978
rect 146678 292294 146734 292350
rect 146802 292294 146858 292350
rect 146678 292170 146734 292226
rect 146802 292170 146858 292226
rect 146678 292046 146734 292102
rect 146802 292046 146858 292102
rect 146678 291922 146734 291978
rect 146802 291922 146858 291978
rect 177398 292294 177454 292350
rect 177522 292294 177578 292350
rect 177398 292170 177454 292226
rect 177522 292170 177578 292226
rect 177398 292046 177454 292102
rect 177522 292046 177578 292102
rect 177398 291922 177454 291978
rect 177522 291922 177578 291978
rect 208118 292294 208174 292350
rect 208242 292294 208298 292350
rect 208118 292170 208174 292226
rect 208242 292170 208298 292226
rect 208118 292046 208174 292102
rect 208242 292046 208298 292102
rect 208118 291922 208174 291978
rect 208242 291922 208298 291978
rect 238838 292294 238894 292350
rect 238962 292294 239018 292350
rect 238838 292170 238894 292226
rect 238962 292170 239018 292226
rect 238838 292046 238894 292102
rect 238962 292046 239018 292102
rect 238838 291922 238894 291978
rect 238962 291922 239018 291978
rect 269558 292294 269614 292350
rect 269682 292294 269738 292350
rect 269558 292170 269614 292226
rect 269682 292170 269738 292226
rect 269558 292046 269614 292102
rect 269682 292046 269738 292102
rect 269558 291922 269614 291978
rect 269682 291922 269738 291978
rect 300278 292294 300334 292350
rect 300402 292294 300458 292350
rect 300278 292170 300334 292226
rect 300402 292170 300458 292226
rect 300278 292046 300334 292102
rect 300402 292046 300458 292102
rect 300278 291922 300334 291978
rect 300402 291922 300458 291978
rect 330998 292294 331054 292350
rect 331122 292294 331178 292350
rect 330998 292170 331054 292226
rect 331122 292170 331178 292226
rect 330998 292046 331054 292102
rect 331122 292046 331178 292102
rect 330998 291922 331054 291978
rect 331122 291922 331178 291978
rect 361718 292294 361774 292350
rect 361842 292294 361898 292350
rect 361718 292170 361774 292226
rect 361842 292170 361898 292226
rect 361718 292046 361774 292102
rect 361842 292046 361898 292102
rect 361718 291922 361774 291978
rect 361842 291922 361898 291978
rect 392438 292294 392494 292350
rect 392562 292294 392618 292350
rect 392438 292170 392494 292226
rect 392562 292170 392618 292226
rect 392438 292046 392494 292102
rect 392562 292046 392618 292102
rect 392438 291922 392494 291978
rect 392562 291922 392618 291978
rect 423158 292294 423214 292350
rect 423282 292294 423338 292350
rect 423158 292170 423214 292226
rect 423282 292170 423338 292226
rect 423158 292046 423214 292102
rect 423282 292046 423338 292102
rect 423158 291922 423214 291978
rect 423282 291922 423338 291978
rect 453878 292294 453934 292350
rect 454002 292294 454058 292350
rect 453878 292170 453934 292226
rect 454002 292170 454058 292226
rect 453878 292046 453934 292102
rect 454002 292046 454058 292102
rect 453878 291922 453934 291978
rect 454002 291922 454058 291978
rect 484598 292294 484654 292350
rect 484722 292294 484778 292350
rect 484598 292170 484654 292226
rect 484722 292170 484778 292226
rect 484598 292046 484654 292102
rect 484722 292046 484778 292102
rect 484598 291922 484654 291978
rect 484722 291922 484778 291978
rect 515318 292294 515374 292350
rect 515442 292294 515498 292350
rect 515318 292170 515374 292226
rect 515442 292170 515498 292226
rect 515318 292046 515374 292102
rect 515442 292046 515498 292102
rect 515318 291922 515374 291978
rect 515442 291922 515498 291978
rect 546038 292294 546094 292350
rect 546162 292294 546218 292350
rect 546038 292170 546094 292226
rect 546162 292170 546218 292226
rect 546038 292046 546094 292102
rect 546162 292046 546218 292102
rect 546038 291922 546094 291978
rect 546162 291922 546218 291978
rect 561250 292294 561306 292350
rect 561374 292294 561430 292350
rect 561498 292294 561554 292350
rect 561622 292294 561678 292350
rect 561250 292170 561306 292226
rect 561374 292170 561430 292226
rect 561498 292170 561554 292226
rect 561622 292170 561678 292226
rect 561250 292046 561306 292102
rect 561374 292046 561430 292102
rect 561498 292046 561554 292102
rect 561622 292046 561678 292102
rect 561250 291922 561306 291978
rect 561374 291922 561430 291978
rect 561498 291922 561554 291978
rect 561622 291922 561678 291978
rect 131318 280294 131374 280350
rect 131442 280294 131498 280350
rect 131318 280170 131374 280226
rect 131442 280170 131498 280226
rect 131318 280046 131374 280102
rect 131442 280046 131498 280102
rect 131318 279922 131374 279978
rect 131442 279922 131498 279978
rect 162038 280294 162094 280350
rect 162162 280294 162218 280350
rect 162038 280170 162094 280226
rect 162162 280170 162218 280226
rect 162038 280046 162094 280102
rect 162162 280046 162218 280102
rect 162038 279922 162094 279978
rect 162162 279922 162218 279978
rect 192758 280294 192814 280350
rect 192882 280294 192938 280350
rect 192758 280170 192814 280226
rect 192882 280170 192938 280226
rect 192758 280046 192814 280102
rect 192882 280046 192938 280102
rect 192758 279922 192814 279978
rect 192882 279922 192938 279978
rect 223478 280294 223534 280350
rect 223602 280294 223658 280350
rect 223478 280170 223534 280226
rect 223602 280170 223658 280226
rect 223478 280046 223534 280102
rect 223602 280046 223658 280102
rect 223478 279922 223534 279978
rect 223602 279922 223658 279978
rect 254198 280294 254254 280350
rect 254322 280294 254378 280350
rect 254198 280170 254254 280226
rect 254322 280170 254378 280226
rect 254198 280046 254254 280102
rect 254322 280046 254378 280102
rect 254198 279922 254254 279978
rect 254322 279922 254378 279978
rect 284918 280294 284974 280350
rect 285042 280294 285098 280350
rect 284918 280170 284974 280226
rect 285042 280170 285098 280226
rect 284918 280046 284974 280102
rect 285042 280046 285098 280102
rect 284918 279922 284974 279978
rect 285042 279922 285098 279978
rect 315638 280294 315694 280350
rect 315762 280294 315818 280350
rect 315638 280170 315694 280226
rect 315762 280170 315818 280226
rect 315638 280046 315694 280102
rect 315762 280046 315818 280102
rect 315638 279922 315694 279978
rect 315762 279922 315818 279978
rect 346358 280294 346414 280350
rect 346482 280294 346538 280350
rect 346358 280170 346414 280226
rect 346482 280170 346538 280226
rect 346358 280046 346414 280102
rect 346482 280046 346538 280102
rect 346358 279922 346414 279978
rect 346482 279922 346538 279978
rect 377078 280294 377134 280350
rect 377202 280294 377258 280350
rect 377078 280170 377134 280226
rect 377202 280170 377258 280226
rect 377078 280046 377134 280102
rect 377202 280046 377258 280102
rect 377078 279922 377134 279978
rect 377202 279922 377258 279978
rect 407798 280294 407854 280350
rect 407922 280294 407978 280350
rect 407798 280170 407854 280226
rect 407922 280170 407978 280226
rect 407798 280046 407854 280102
rect 407922 280046 407978 280102
rect 407798 279922 407854 279978
rect 407922 279922 407978 279978
rect 438518 280294 438574 280350
rect 438642 280294 438698 280350
rect 438518 280170 438574 280226
rect 438642 280170 438698 280226
rect 438518 280046 438574 280102
rect 438642 280046 438698 280102
rect 438518 279922 438574 279978
rect 438642 279922 438698 279978
rect 469238 280294 469294 280350
rect 469362 280294 469418 280350
rect 469238 280170 469294 280226
rect 469362 280170 469418 280226
rect 469238 280046 469294 280102
rect 469362 280046 469418 280102
rect 469238 279922 469294 279978
rect 469362 279922 469418 279978
rect 499958 280294 500014 280350
rect 500082 280294 500138 280350
rect 499958 280170 500014 280226
rect 500082 280170 500138 280226
rect 499958 280046 500014 280102
rect 500082 280046 500138 280102
rect 499958 279922 500014 279978
rect 500082 279922 500138 279978
rect 530678 280294 530734 280350
rect 530802 280294 530858 280350
rect 530678 280170 530734 280226
rect 530802 280170 530858 280226
rect 530678 280046 530734 280102
rect 530802 280046 530858 280102
rect 530678 279922 530734 279978
rect 530802 279922 530858 279978
rect 111250 274294 111306 274350
rect 111374 274294 111430 274350
rect 111498 274294 111554 274350
rect 111622 274294 111678 274350
rect 111250 274170 111306 274226
rect 111374 274170 111430 274226
rect 111498 274170 111554 274226
rect 111622 274170 111678 274226
rect 111250 274046 111306 274102
rect 111374 274046 111430 274102
rect 111498 274046 111554 274102
rect 111622 274046 111678 274102
rect 111250 273922 111306 273978
rect 111374 273922 111430 273978
rect 111498 273922 111554 273978
rect 111622 273922 111678 273978
rect 96970 262294 97026 262350
rect 97094 262294 97150 262350
rect 97218 262294 97274 262350
rect 97342 262294 97398 262350
rect 96970 262170 97026 262226
rect 97094 262170 97150 262226
rect 97218 262170 97274 262226
rect 97342 262170 97398 262226
rect 96970 262046 97026 262102
rect 97094 262046 97150 262102
rect 97218 262046 97274 262102
rect 97342 262046 97398 262102
rect 96970 261922 97026 261978
rect 97094 261922 97150 261978
rect 97218 261922 97274 261978
rect 97342 261922 97398 261978
rect 100598 262294 100654 262350
rect 100722 262294 100778 262350
rect 100598 262170 100654 262226
rect 100722 262170 100778 262226
rect 100598 262046 100654 262102
rect 100722 262046 100778 262102
rect 100598 261922 100654 261978
rect 100722 261922 100778 261978
rect 115958 274294 116014 274350
rect 116082 274294 116138 274350
rect 115958 274170 116014 274226
rect 116082 274170 116138 274226
rect 115958 274046 116014 274102
rect 116082 274046 116138 274102
rect 115958 273922 116014 273978
rect 116082 273922 116138 273978
rect 146678 274294 146734 274350
rect 146802 274294 146858 274350
rect 146678 274170 146734 274226
rect 146802 274170 146858 274226
rect 146678 274046 146734 274102
rect 146802 274046 146858 274102
rect 146678 273922 146734 273978
rect 146802 273922 146858 273978
rect 177398 274294 177454 274350
rect 177522 274294 177578 274350
rect 177398 274170 177454 274226
rect 177522 274170 177578 274226
rect 177398 274046 177454 274102
rect 177522 274046 177578 274102
rect 177398 273922 177454 273978
rect 177522 273922 177578 273978
rect 208118 274294 208174 274350
rect 208242 274294 208298 274350
rect 208118 274170 208174 274226
rect 208242 274170 208298 274226
rect 208118 274046 208174 274102
rect 208242 274046 208298 274102
rect 208118 273922 208174 273978
rect 208242 273922 208298 273978
rect 238838 274294 238894 274350
rect 238962 274294 239018 274350
rect 238838 274170 238894 274226
rect 238962 274170 239018 274226
rect 238838 274046 238894 274102
rect 238962 274046 239018 274102
rect 238838 273922 238894 273978
rect 238962 273922 239018 273978
rect 269558 274294 269614 274350
rect 269682 274294 269738 274350
rect 269558 274170 269614 274226
rect 269682 274170 269738 274226
rect 269558 274046 269614 274102
rect 269682 274046 269738 274102
rect 269558 273922 269614 273978
rect 269682 273922 269738 273978
rect 300278 274294 300334 274350
rect 300402 274294 300458 274350
rect 300278 274170 300334 274226
rect 300402 274170 300458 274226
rect 300278 274046 300334 274102
rect 300402 274046 300458 274102
rect 300278 273922 300334 273978
rect 300402 273922 300458 273978
rect 330998 274294 331054 274350
rect 331122 274294 331178 274350
rect 330998 274170 331054 274226
rect 331122 274170 331178 274226
rect 330998 274046 331054 274102
rect 331122 274046 331178 274102
rect 330998 273922 331054 273978
rect 331122 273922 331178 273978
rect 361718 274294 361774 274350
rect 361842 274294 361898 274350
rect 361718 274170 361774 274226
rect 361842 274170 361898 274226
rect 361718 274046 361774 274102
rect 361842 274046 361898 274102
rect 361718 273922 361774 273978
rect 361842 273922 361898 273978
rect 392438 274294 392494 274350
rect 392562 274294 392618 274350
rect 392438 274170 392494 274226
rect 392562 274170 392618 274226
rect 392438 274046 392494 274102
rect 392562 274046 392618 274102
rect 392438 273922 392494 273978
rect 392562 273922 392618 273978
rect 423158 274294 423214 274350
rect 423282 274294 423338 274350
rect 423158 274170 423214 274226
rect 423282 274170 423338 274226
rect 423158 274046 423214 274102
rect 423282 274046 423338 274102
rect 423158 273922 423214 273978
rect 423282 273922 423338 273978
rect 453878 274294 453934 274350
rect 454002 274294 454058 274350
rect 453878 274170 453934 274226
rect 454002 274170 454058 274226
rect 453878 274046 453934 274102
rect 454002 274046 454058 274102
rect 453878 273922 453934 273978
rect 454002 273922 454058 273978
rect 484598 274294 484654 274350
rect 484722 274294 484778 274350
rect 484598 274170 484654 274226
rect 484722 274170 484778 274226
rect 484598 274046 484654 274102
rect 484722 274046 484778 274102
rect 484598 273922 484654 273978
rect 484722 273922 484778 273978
rect 515318 274294 515374 274350
rect 515442 274294 515498 274350
rect 515318 274170 515374 274226
rect 515442 274170 515498 274226
rect 515318 274046 515374 274102
rect 515442 274046 515498 274102
rect 515318 273922 515374 273978
rect 515442 273922 515498 273978
rect 546038 274294 546094 274350
rect 546162 274294 546218 274350
rect 546038 274170 546094 274226
rect 546162 274170 546218 274226
rect 546038 274046 546094 274102
rect 546162 274046 546218 274102
rect 546038 273922 546094 273978
rect 546162 273922 546218 273978
rect 561250 274294 561306 274350
rect 561374 274294 561430 274350
rect 561498 274294 561554 274350
rect 561622 274294 561678 274350
rect 561250 274170 561306 274226
rect 561374 274170 561430 274226
rect 561498 274170 561554 274226
rect 561622 274170 561678 274226
rect 561250 274046 561306 274102
rect 561374 274046 561430 274102
rect 561498 274046 561554 274102
rect 561622 274046 561678 274102
rect 561250 273922 561306 273978
rect 561374 273922 561430 273978
rect 561498 273922 561554 273978
rect 561622 273922 561678 273978
rect 131318 262294 131374 262350
rect 131442 262294 131498 262350
rect 131318 262170 131374 262226
rect 131442 262170 131498 262226
rect 131318 262046 131374 262102
rect 131442 262046 131498 262102
rect 131318 261922 131374 261978
rect 131442 261922 131498 261978
rect 162038 262294 162094 262350
rect 162162 262294 162218 262350
rect 162038 262170 162094 262226
rect 162162 262170 162218 262226
rect 162038 262046 162094 262102
rect 162162 262046 162218 262102
rect 162038 261922 162094 261978
rect 162162 261922 162218 261978
rect 192758 262294 192814 262350
rect 192882 262294 192938 262350
rect 192758 262170 192814 262226
rect 192882 262170 192938 262226
rect 192758 262046 192814 262102
rect 192882 262046 192938 262102
rect 192758 261922 192814 261978
rect 192882 261922 192938 261978
rect 223478 262294 223534 262350
rect 223602 262294 223658 262350
rect 223478 262170 223534 262226
rect 223602 262170 223658 262226
rect 223478 262046 223534 262102
rect 223602 262046 223658 262102
rect 223478 261922 223534 261978
rect 223602 261922 223658 261978
rect 254198 262294 254254 262350
rect 254322 262294 254378 262350
rect 254198 262170 254254 262226
rect 254322 262170 254378 262226
rect 254198 262046 254254 262102
rect 254322 262046 254378 262102
rect 254198 261922 254254 261978
rect 254322 261922 254378 261978
rect 284918 262294 284974 262350
rect 285042 262294 285098 262350
rect 284918 262170 284974 262226
rect 285042 262170 285098 262226
rect 284918 262046 284974 262102
rect 285042 262046 285098 262102
rect 284918 261922 284974 261978
rect 285042 261922 285098 261978
rect 315638 262294 315694 262350
rect 315762 262294 315818 262350
rect 315638 262170 315694 262226
rect 315762 262170 315818 262226
rect 315638 262046 315694 262102
rect 315762 262046 315818 262102
rect 315638 261922 315694 261978
rect 315762 261922 315818 261978
rect 346358 262294 346414 262350
rect 346482 262294 346538 262350
rect 346358 262170 346414 262226
rect 346482 262170 346538 262226
rect 346358 262046 346414 262102
rect 346482 262046 346538 262102
rect 346358 261922 346414 261978
rect 346482 261922 346538 261978
rect 377078 262294 377134 262350
rect 377202 262294 377258 262350
rect 377078 262170 377134 262226
rect 377202 262170 377258 262226
rect 377078 262046 377134 262102
rect 377202 262046 377258 262102
rect 377078 261922 377134 261978
rect 377202 261922 377258 261978
rect 407798 262294 407854 262350
rect 407922 262294 407978 262350
rect 407798 262170 407854 262226
rect 407922 262170 407978 262226
rect 407798 262046 407854 262102
rect 407922 262046 407978 262102
rect 407798 261922 407854 261978
rect 407922 261922 407978 261978
rect 438518 262294 438574 262350
rect 438642 262294 438698 262350
rect 438518 262170 438574 262226
rect 438642 262170 438698 262226
rect 438518 262046 438574 262102
rect 438642 262046 438698 262102
rect 438518 261922 438574 261978
rect 438642 261922 438698 261978
rect 469238 262294 469294 262350
rect 469362 262294 469418 262350
rect 469238 262170 469294 262226
rect 469362 262170 469418 262226
rect 469238 262046 469294 262102
rect 469362 262046 469418 262102
rect 469238 261922 469294 261978
rect 469362 261922 469418 261978
rect 499958 262294 500014 262350
rect 500082 262294 500138 262350
rect 499958 262170 500014 262226
rect 500082 262170 500138 262226
rect 499958 262046 500014 262102
rect 500082 262046 500138 262102
rect 499958 261922 500014 261978
rect 500082 261922 500138 261978
rect 530678 262294 530734 262350
rect 530802 262294 530858 262350
rect 530678 262170 530734 262226
rect 530802 262170 530858 262226
rect 530678 262046 530734 262102
rect 530802 262046 530858 262102
rect 530678 261922 530734 261978
rect 530802 261922 530858 261978
rect 111250 256294 111306 256350
rect 111374 256294 111430 256350
rect 111498 256294 111554 256350
rect 111622 256294 111678 256350
rect 111250 256170 111306 256226
rect 111374 256170 111430 256226
rect 111498 256170 111554 256226
rect 111622 256170 111678 256226
rect 111250 256046 111306 256102
rect 111374 256046 111430 256102
rect 111498 256046 111554 256102
rect 111622 256046 111678 256102
rect 111250 255922 111306 255978
rect 111374 255922 111430 255978
rect 111498 255922 111554 255978
rect 111622 255922 111678 255978
rect 96970 244294 97026 244350
rect 97094 244294 97150 244350
rect 97218 244294 97274 244350
rect 97342 244294 97398 244350
rect 96970 244170 97026 244226
rect 97094 244170 97150 244226
rect 97218 244170 97274 244226
rect 97342 244170 97398 244226
rect 96970 244046 97026 244102
rect 97094 244046 97150 244102
rect 97218 244046 97274 244102
rect 97342 244046 97398 244102
rect 96970 243922 97026 243978
rect 97094 243922 97150 243978
rect 97218 243922 97274 243978
rect 97342 243922 97398 243978
rect 100598 244294 100654 244350
rect 100722 244294 100778 244350
rect 100598 244170 100654 244226
rect 100722 244170 100778 244226
rect 100598 244046 100654 244102
rect 100722 244046 100778 244102
rect 100598 243922 100654 243978
rect 100722 243922 100778 243978
rect 115958 256294 116014 256350
rect 116082 256294 116138 256350
rect 115958 256170 116014 256226
rect 116082 256170 116138 256226
rect 115958 256046 116014 256102
rect 116082 256046 116138 256102
rect 115958 255922 116014 255978
rect 116082 255922 116138 255978
rect 146678 256294 146734 256350
rect 146802 256294 146858 256350
rect 146678 256170 146734 256226
rect 146802 256170 146858 256226
rect 146678 256046 146734 256102
rect 146802 256046 146858 256102
rect 146678 255922 146734 255978
rect 146802 255922 146858 255978
rect 177398 256294 177454 256350
rect 177522 256294 177578 256350
rect 177398 256170 177454 256226
rect 177522 256170 177578 256226
rect 177398 256046 177454 256102
rect 177522 256046 177578 256102
rect 177398 255922 177454 255978
rect 177522 255922 177578 255978
rect 208118 256294 208174 256350
rect 208242 256294 208298 256350
rect 208118 256170 208174 256226
rect 208242 256170 208298 256226
rect 208118 256046 208174 256102
rect 208242 256046 208298 256102
rect 208118 255922 208174 255978
rect 208242 255922 208298 255978
rect 238838 256294 238894 256350
rect 238962 256294 239018 256350
rect 238838 256170 238894 256226
rect 238962 256170 239018 256226
rect 238838 256046 238894 256102
rect 238962 256046 239018 256102
rect 238838 255922 238894 255978
rect 238962 255922 239018 255978
rect 269558 256294 269614 256350
rect 269682 256294 269738 256350
rect 269558 256170 269614 256226
rect 269682 256170 269738 256226
rect 269558 256046 269614 256102
rect 269682 256046 269738 256102
rect 269558 255922 269614 255978
rect 269682 255922 269738 255978
rect 300278 256294 300334 256350
rect 300402 256294 300458 256350
rect 300278 256170 300334 256226
rect 300402 256170 300458 256226
rect 300278 256046 300334 256102
rect 300402 256046 300458 256102
rect 300278 255922 300334 255978
rect 300402 255922 300458 255978
rect 330998 256294 331054 256350
rect 331122 256294 331178 256350
rect 330998 256170 331054 256226
rect 331122 256170 331178 256226
rect 330998 256046 331054 256102
rect 331122 256046 331178 256102
rect 330998 255922 331054 255978
rect 331122 255922 331178 255978
rect 361718 256294 361774 256350
rect 361842 256294 361898 256350
rect 361718 256170 361774 256226
rect 361842 256170 361898 256226
rect 361718 256046 361774 256102
rect 361842 256046 361898 256102
rect 361718 255922 361774 255978
rect 361842 255922 361898 255978
rect 392438 256294 392494 256350
rect 392562 256294 392618 256350
rect 392438 256170 392494 256226
rect 392562 256170 392618 256226
rect 392438 256046 392494 256102
rect 392562 256046 392618 256102
rect 392438 255922 392494 255978
rect 392562 255922 392618 255978
rect 423158 256294 423214 256350
rect 423282 256294 423338 256350
rect 423158 256170 423214 256226
rect 423282 256170 423338 256226
rect 423158 256046 423214 256102
rect 423282 256046 423338 256102
rect 423158 255922 423214 255978
rect 423282 255922 423338 255978
rect 453878 256294 453934 256350
rect 454002 256294 454058 256350
rect 453878 256170 453934 256226
rect 454002 256170 454058 256226
rect 453878 256046 453934 256102
rect 454002 256046 454058 256102
rect 453878 255922 453934 255978
rect 454002 255922 454058 255978
rect 484598 256294 484654 256350
rect 484722 256294 484778 256350
rect 484598 256170 484654 256226
rect 484722 256170 484778 256226
rect 484598 256046 484654 256102
rect 484722 256046 484778 256102
rect 484598 255922 484654 255978
rect 484722 255922 484778 255978
rect 515318 256294 515374 256350
rect 515442 256294 515498 256350
rect 515318 256170 515374 256226
rect 515442 256170 515498 256226
rect 515318 256046 515374 256102
rect 515442 256046 515498 256102
rect 515318 255922 515374 255978
rect 515442 255922 515498 255978
rect 546038 256294 546094 256350
rect 546162 256294 546218 256350
rect 546038 256170 546094 256226
rect 546162 256170 546218 256226
rect 546038 256046 546094 256102
rect 546162 256046 546218 256102
rect 546038 255922 546094 255978
rect 546162 255922 546218 255978
rect 561250 256294 561306 256350
rect 561374 256294 561430 256350
rect 561498 256294 561554 256350
rect 561622 256294 561678 256350
rect 561250 256170 561306 256226
rect 561374 256170 561430 256226
rect 561498 256170 561554 256226
rect 561622 256170 561678 256226
rect 561250 256046 561306 256102
rect 561374 256046 561430 256102
rect 561498 256046 561554 256102
rect 561622 256046 561678 256102
rect 561250 255922 561306 255978
rect 561374 255922 561430 255978
rect 561498 255922 561554 255978
rect 561622 255922 561678 255978
rect 131318 244294 131374 244350
rect 131442 244294 131498 244350
rect 131318 244170 131374 244226
rect 131442 244170 131498 244226
rect 131318 244046 131374 244102
rect 131442 244046 131498 244102
rect 131318 243922 131374 243978
rect 131442 243922 131498 243978
rect 162038 244294 162094 244350
rect 162162 244294 162218 244350
rect 162038 244170 162094 244226
rect 162162 244170 162218 244226
rect 162038 244046 162094 244102
rect 162162 244046 162218 244102
rect 162038 243922 162094 243978
rect 162162 243922 162218 243978
rect 192758 244294 192814 244350
rect 192882 244294 192938 244350
rect 192758 244170 192814 244226
rect 192882 244170 192938 244226
rect 192758 244046 192814 244102
rect 192882 244046 192938 244102
rect 192758 243922 192814 243978
rect 192882 243922 192938 243978
rect 223478 244294 223534 244350
rect 223602 244294 223658 244350
rect 223478 244170 223534 244226
rect 223602 244170 223658 244226
rect 223478 244046 223534 244102
rect 223602 244046 223658 244102
rect 223478 243922 223534 243978
rect 223602 243922 223658 243978
rect 254198 244294 254254 244350
rect 254322 244294 254378 244350
rect 254198 244170 254254 244226
rect 254322 244170 254378 244226
rect 254198 244046 254254 244102
rect 254322 244046 254378 244102
rect 254198 243922 254254 243978
rect 254322 243922 254378 243978
rect 284918 244294 284974 244350
rect 285042 244294 285098 244350
rect 284918 244170 284974 244226
rect 285042 244170 285098 244226
rect 284918 244046 284974 244102
rect 285042 244046 285098 244102
rect 284918 243922 284974 243978
rect 285042 243922 285098 243978
rect 315638 244294 315694 244350
rect 315762 244294 315818 244350
rect 315638 244170 315694 244226
rect 315762 244170 315818 244226
rect 315638 244046 315694 244102
rect 315762 244046 315818 244102
rect 315638 243922 315694 243978
rect 315762 243922 315818 243978
rect 346358 244294 346414 244350
rect 346482 244294 346538 244350
rect 346358 244170 346414 244226
rect 346482 244170 346538 244226
rect 346358 244046 346414 244102
rect 346482 244046 346538 244102
rect 346358 243922 346414 243978
rect 346482 243922 346538 243978
rect 377078 244294 377134 244350
rect 377202 244294 377258 244350
rect 377078 244170 377134 244226
rect 377202 244170 377258 244226
rect 377078 244046 377134 244102
rect 377202 244046 377258 244102
rect 377078 243922 377134 243978
rect 377202 243922 377258 243978
rect 407798 244294 407854 244350
rect 407922 244294 407978 244350
rect 407798 244170 407854 244226
rect 407922 244170 407978 244226
rect 407798 244046 407854 244102
rect 407922 244046 407978 244102
rect 407798 243922 407854 243978
rect 407922 243922 407978 243978
rect 438518 244294 438574 244350
rect 438642 244294 438698 244350
rect 438518 244170 438574 244226
rect 438642 244170 438698 244226
rect 438518 244046 438574 244102
rect 438642 244046 438698 244102
rect 438518 243922 438574 243978
rect 438642 243922 438698 243978
rect 469238 244294 469294 244350
rect 469362 244294 469418 244350
rect 469238 244170 469294 244226
rect 469362 244170 469418 244226
rect 469238 244046 469294 244102
rect 469362 244046 469418 244102
rect 469238 243922 469294 243978
rect 469362 243922 469418 243978
rect 499958 244294 500014 244350
rect 500082 244294 500138 244350
rect 499958 244170 500014 244226
rect 500082 244170 500138 244226
rect 499958 244046 500014 244102
rect 500082 244046 500138 244102
rect 499958 243922 500014 243978
rect 500082 243922 500138 243978
rect 530678 244294 530734 244350
rect 530802 244294 530858 244350
rect 530678 244170 530734 244226
rect 530802 244170 530858 244226
rect 530678 244046 530734 244102
rect 530802 244046 530858 244102
rect 530678 243922 530734 243978
rect 530802 243922 530858 243978
rect 111250 238294 111306 238350
rect 111374 238294 111430 238350
rect 111498 238294 111554 238350
rect 111622 238294 111678 238350
rect 111250 238170 111306 238226
rect 111374 238170 111430 238226
rect 111498 238170 111554 238226
rect 111622 238170 111678 238226
rect 111250 238046 111306 238102
rect 111374 238046 111430 238102
rect 111498 238046 111554 238102
rect 111622 238046 111678 238102
rect 111250 237922 111306 237978
rect 111374 237922 111430 237978
rect 111498 237922 111554 237978
rect 111622 237922 111678 237978
rect 96970 226294 97026 226350
rect 97094 226294 97150 226350
rect 97218 226294 97274 226350
rect 97342 226294 97398 226350
rect 96970 226170 97026 226226
rect 97094 226170 97150 226226
rect 97218 226170 97274 226226
rect 97342 226170 97398 226226
rect 96970 226046 97026 226102
rect 97094 226046 97150 226102
rect 97218 226046 97274 226102
rect 97342 226046 97398 226102
rect 96970 225922 97026 225978
rect 97094 225922 97150 225978
rect 97218 225922 97274 225978
rect 97342 225922 97398 225978
rect 100598 226294 100654 226350
rect 100722 226294 100778 226350
rect 100598 226170 100654 226226
rect 100722 226170 100778 226226
rect 100598 226046 100654 226102
rect 100722 226046 100778 226102
rect 100598 225922 100654 225978
rect 100722 225922 100778 225978
rect 115958 238294 116014 238350
rect 116082 238294 116138 238350
rect 115958 238170 116014 238226
rect 116082 238170 116138 238226
rect 115958 238046 116014 238102
rect 116082 238046 116138 238102
rect 115958 237922 116014 237978
rect 116082 237922 116138 237978
rect 146678 238294 146734 238350
rect 146802 238294 146858 238350
rect 146678 238170 146734 238226
rect 146802 238170 146858 238226
rect 146678 238046 146734 238102
rect 146802 238046 146858 238102
rect 146678 237922 146734 237978
rect 146802 237922 146858 237978
rect 177398 238294 177454 238350
rect 177522 238294 177578 238350
rect 177398 238170 177454 238226
rect 177522 238170 177578 238226
rect 177398 238046 177454 238102
rect 177522 238046 177578 238102
rect 177398 237922 177454 237978
rect 177522 237922 177578 237978
rect 208118 238294 208174 238350
rect 208242 238294 208298 238350
rect 208118 238170 208174 238226
rect 208242 238170 208298 238226
rect 208118 238046 208174 238102
rect 208242 238046 208298 238102
rect 208118 237922 208174 237978
rect 208242 237922 208298 237978
rect 238838 238294 238894 238350
rect 238962 238294 239018 238350
rect 238838 238170 238894 238226
rect 238962 238170 239018 238226
rect 238838 238046 238894 238102
rect 238962 238046 239018 238102
rect 238838 237922 238894 237978
rect 238962 237922 239018 237978
rect 269558 238294 269614 238350
rect 269682 238294 269738 238350
rect 269558 238170 269614 238226
rect 269682 238170 269738 238226
rect 269558 238046 269614 238102
rect 269682 238046 269738 238102
rect 269558 237922 269614 237978
rect 269682 237922 269738 237978
rect 300278 238294 300334 238350
rect 300402 238294 300458 238350
rect 300278 238170 300334 238226
rect 300402 238170 300458 238226
rect 300278 238046 300334 238102
rect 300402 238046 300458 238102
rect 300278 237922 300334 237978
rect 300402 237922 300458 237978
rect 330998 238294 331054 238350
rect 331122 238294 331178 238350
rect 330998 238170 331054 238226
rect 331122 238170 331178 238226
rect 330998 238046 331054 238102
rect 331122 238046 331178 238102
rect 330998 237922 331054 237978
rect 331122 237922 331178 237978
rect 361718 238294 361774 238350
rect 361842 238294 361898 238350
rect 361718 238170 361774 238226
rect 361842 238170 361898 238226
rect 361718 238046 361774 238102
rect 361842 238046 361898 238102
rect 361718 237922 361774 237978
rect 361842 237922 361898 237978
rect 392438 238294 392494 238350
rect 392562 238294 392618 238350
rect 392438 238170 392494 238226
rect 392562 238170 392618 238226
rect 392438 238046 392494 238102
rect 392562 238046 392618 238102
rect 392438 237922 392494 237978
rect 392562 237922 392618 237978
rect 423158 238294 423214 238350
rect 423282 238294 423338 238350
rect 423158 238170 423214 238226
rect 423282 238170 423338 238226
rect 423158 238046 423214 238102
rect 423282 238046 423338 238102
rect 423158 237922 423214 237978
rect 423282 237922 423338 237978
rect 453878 238294 453934 238350
rect 454002 238294 454058 238350
rect 453878 238170 453934 238226
rect 454002 238170 454058 238226
rect 453878 238046 453934 238102
rect 454002 238046 454058 238102
rect 453878 237922 453934 237978
rect 454002 237922 454058 237978
rect 484598 238294 484654 238350
rect 484722 238294 484778 238350
rect 484598 238170 484654 238226
rect 484722 238170 484778 238226
rect 484598 238046 484654 238102
rect 484722 238046 484778 238102
rect 484598 237922 484654 237978
rect 484722 237922 484778 237978
rect 515318 238294 515374 238350
rect 515442 238294 515498 238350
rect 515318 238170 515374 238226
rect 515442 238170 515498 238226
rect 515318 238046 515374 238102
rect 515442 238046 515498 238102
rect 515318 237922 515374 237978
rect 515442 237922 515498 237978
rect 546038 238294 546094 238350
rect 546162 238294 546218 238350
rect 546038 238170 546094 238226
rect 546162 238170 546218 238226
rect 546038 238046 546094 238102
rect 546162 238046 546218 238102
rect 546038 237922 546094 237978
rect 546162 237922 546218 237978
rect 561250 238294 561306 238350
rect 561374 238294 561430 238350
rect 561498 238294 561554 238350
rect 561622 238294 561678 238350
rect 561250 238170 561306 238226
rect 561374 238170 561430 238226
rect 561498 238170 561554 238226
rect 561622 238170 561678 238226
rect 561250 238046 561306 238102
rect 561374 238046 561430 238102
rect 561498 238046 561554 238102
rect 561622 238046 561678 238102
rect 561250 237922 561306 237978
rect 561374 237922 561430 237978
rect 561498 237922 561554 237978
rect 561622 237922 561678 237978
rect 131318 226294 131374 226350
rect 131442 226294 131498 226350
rect 131318 226170 131374 226226
rect 131442 226170 131498 226226
rect 131318 226046 131374 226102
rect 131442 226046 131498 226102
rect 131318 225922 131374 225978
rect 131442 225922 131498 225978
rect 162038 226294 162094 226350
rect 162162 226294 162218 226350
rect 162038 226170 162094 226226
rect 162162 226170 162218 226226
rect 162038 226046 162094 226102
rect 162162 226046 162218 226102
rect 162038 225922 162094 225978
rect 162162 225922 162218 225978
rect 192758 226294 192814 226350
rect 192882 226294 192938 226350
rect 192758 226170 192814 226226
rect 192882 226170 192938 226226
rect 192758 226046 192814 226102
rect 192882 226046 192938 226102
rect 192758 225922 192814 225978
rect 192882 225922 192938 225978
rect 223478 226294 223534 226350
rect 223602 226294 223658 226350
rect 223478 226170 223534 226226
rect 223602 226170 223658 226226
rect 223478 226046 223534 226102
rect 223602 226046 223658 226102
rect 223478 225922 223534 225978
rect 223602 225922 223658 225978
rect 254198 226294 254254 226350
rect 254322 226294 254378 226350
rect 254198 226170 254254 226226
rect 254322 226170 254378 226226
rect 254198 226046 254254 226102
rect 254322 226046 254378 226102
rect 254198 225922 254254 225978
rect 254322 225922 254378 225978
rect 284918 226294 284974 226350
rect 285042 226294 285098 226350
rect 284918 226170 284974 226226
rect 285042 226170 285098 226226
rect 284918 226046 284974 226102
rect 285042 226046 285098 226102
rect 284918 225922 284974 225978
rect 285042 225922 285098 225978
rect 315638 226294 315694 226350
rect 315762 226294 315818 226350
rect 315638 226170 315694 226226
rect 315762 226170 315818 226226
rect 315638 226046 315694 226102
rect 315762 226046 315818 226102
rect 315638 225922 315694 225978
rect 315762 225922 315818 225978
rect 346358 226294 346414 226350
rect 346482 226294 346538 226350
rect 346358 226170 346414 226226
rect 346482 226170 346538 226226
rect 346358 226046 346414 226102
rect 346482 226046 346538 226102
rect 346358 225922 346414 225978
rect 346482 225922 346538 225978
rect 377078 226294 377134 226350
rect 377202 226294 377258 226350
rect 377078 226170 377134 226226
rect 377202 226170 377258 226226
rect 377078 226046 377134 226102
rect 377202 226046 377258 226102
rect 377078 225922 377134 225978
rect 377202 225922 377258 225978
rect 407798 226294 407854 226350
rect 407922 226294 407978 226350
rect 407798 226170 407854 226226
rect 407922 226170 407978 226226
rect 407798 226046 407854 226102
rect 407922 226046 407978 226102
rect 407798 225922 407854 225978
rect 407922 225922 407978 225978
rect 438518 226294 438574 226350
rect 438642 226294 438698 226350
rect 438518 226170 438574 226226
rect 438642 226170 438698 226226
rect 438518 226046 438574 226102
rect 438642 226046 438698 226102
rect 438518 225922 438574 225978
rect 438642 225922 438698 225978
rect 469238 226294 469294 226350
rect 469362 226294 469418 226350
rect 469238 226170 469294 226226
rect 469362 226170 469418 226226
rect 469238 226046 469294 226102
rect 469362 226046 469418 226102
rect 469238 225922 469294 225978
rect 469362 225922 469418 225978
rect 499958 226294 500014 226350
rect 500082 226294 500138 226350
rect 499958 226170 500014 226226
rect 500082 226170 500138 226226
rect 499958 226046 500014 226102
rect 500082 226046 500138 226102
rect 499958 225922 500014 225978
rect 500082 225922 500138 225978
rect 530678 226294 530734 226350
rect 530802 226294 530858 226350
rect 530678 226170 530734 226226
rect 530802 226170 530858 226226
rect 530678 226046 530734 226102
rect 530802 226046 530858 226102
rect 530678 225922 530734 225978
rect 530802 225922 530858 225978
rect 111250 220294 111306 220350
rect 111374 220294 111430 220350
rect 111498 220294 111554 220350
rect 111622 220294 111678 220350
rect 111250 220170 111306 220226
rect 111374 220170 111430 220226
rect 111498 220170 111554 220226
rect 111622 220170 111678 220226
rect 111250 220046 111306 220102
rect 111374 220046 111430 220102
rect 111498 220046 111554 220102
rect 111622 220046 111678 220102
rect 111250 219922 111306 219978
rect 111374 219922 111430 219978
rect 111498 219922 111554 219978
rect 111622 219922 111678 219978
rect 96970 208294 97026 208350
rect 97094 208294 97150 208350
rect 97218 208294 97274 208350
rect 97342 208294 97398 208350
rect 96970 208170 97026 208226
rect 97094 208170 97150 208226
rect 97218 208170 97274 208226
rect 97342 208170 97398 208226
rect 96970 208046 97026 208102
rect 97094 208046 97150 208102
rect 97218 208046 97274 208102
rect 97342 208046 97398 208102
rect 96970 207922 97026 207978
rect 97094 207922 97150 207978
rect 97218 207922 97274 207978
rect 97342 207922 97398 207978
rect 100598 208294 100654 208350
rect 100722 208294 100778 208350
rect 100598 208170 100654 208226
rect 100722 208170 100778 208226
rect 100598 208046 100654 208102
rect 100722 208046 100778 208102
rect 100598 207922 100654 207978
rect 100722 207922 100778 207978
rect 115958 220294 116014 220350
rect 116082 220294 116138 220350
rect 115958 220170 116014 220226
rect 116082 220170 116138 220226
rect 115958 220046 116014 220102
rect 116082 220046 116138 220102
rect 115958 219922 116014 219978
rect 116082 219922 116138 219978
rect 146678 220294 146734 220350
rect 146802 220294 146858 220350
rect 146678 220170 146734 220226
rect 146802 220170 146858 220226
rect 146678 220046 146734 220102
rect 146802 220046 146858 220102
rect 146678 219922 146734 219978
rect 146802 219922 146858 219978
rect 177398 220294 177454 220350
rect 177522 220294 177578 220350
rect 177398 220170 177454 220226
rect 177522 220170 177578 220226
rect 177398 220046 177454 220102
rect 177522 220046 177578 220102
rect 177398 219922 177454 219978
rect 177522 219922 177578 219978
rect 208118 220294 208174 220350
rect 208242 220294 208298 220350
rect 208118 220170 208174 220226
rect 208242 220170 208298 220226
rect 208118 220046 208174 220102
rect 208242 220046 208298 220102
rect 208118 219922 208174 219978
rect 208242 219922 208298 219978
rect 238838 220294 238894 220350
rect 238962 220294 239018 220350
rect 238838 220170 238894 220226
rect 238962 220170 239018 220226
rect 238838 220046 238894 220102
rect 238962 220046 239018 220102
rect 238838 219922 238894 219978
rect 238962 219922 239018 219978
rect 269558 220294 269614 220350
rect 269682 220294 269738 220350
rect 269558 220170 269614 220226
rect 269682 220170 269738 220226
rect 269558 220046 269614 220102
rect 269682 220046 269738 220102
rect 269558 219922 269614 219978
rect 269682 219922 269738 219978
rect 300278 220294 300334 220350
rect 300402 220294 300458 220350
rect 300278 220170 300334 220226
rect 300402 220170 300458 220226
rect 300278 220046 300334 220102
rect 300402 220046 300458 220102
rect 300278 219922 300334 219978
rect 300402 219922 300458 219978
rect 330998 220294 331054 220350
rect 331122 220294 331178 220350
rect 330998 220170 331054 220226
rect 331122 220170 331178 220226
rect 330998 220046 331054 220102
rect 331122 220046 331178 220102
rect 330998 219922 331054 219978
rect 331122 219922 331178 219978
rect 361718 220294 361774 220350
rect 361842 220294 361898 220350
rect 361718 220170 361774 220226
rect 361842 220170 361898 220226
rect 361718 220046 361774 220102
rect 361842 220046 361898 220102
rect 361718 219922 361774 219978
rect 361842 219922 361898 219978
rect 392438 220294 392494 220350
rect 392562 220294 392618 220350
rect 392438 220170 392494 220226
rect 392562 220170 392618 220226
rect 392438 220046 392494 220102
rect 392562 220046 392618 220102
rect 392438 219922 392494 219978
rect 392562 219922 392618 219978
rect 423158 220294 423214 220350
rect 423282 220294 423338 220350
rect 423158 220170 423214 220226
rect 423282 220170 423338 220226
rect 423158 220046 423214 220102
rect 423282 220046 423338 220102
rect 423158 219922 423214 219978
rect 423282 219922 423338 219978
rect 453878 220294 453934 220350
rect 454002 220294 454058 220350
rect 453878 220170 453934 220226
rect 454002 220170 454058 220226
rect 453878 220046 453934 220102
rect 454002 220046 454058 220102
rect 453878 219922 453934 219978
rect 454002 219922 454058 219978
rect 484598 220294 484654 220350
rect 484722 220294 484778 220350
rect 484598 220170 484654 220226
rect 484722 220170 484778 220226
rect 484598 220046 484654 220102
rect 484722 220046 484778 220102
rect 484598 219922 484654 219978
rect 484722 219922 484778 219978
rect 515318 220294 515374 220350
rect 515442 220294 515498 220350
rect 515318 220170 515374 220226
rect 515442 220170 515498 220226
rect 515318 220046 515374 220102
rect 515442 220046 515498 220102
rect 515318 219922 515374 219978
rect 515442 219922 515498 219978
rect 546038 220294 546094 220350
rect 546162 220294 546218 220350
rect 546038 220170 546094 220226
rect 546162 220170 546218 220226
rect 546038 220046 546094 220102
rect 546162 220046 546218 220102
rect 546038 219922 546094 219978
rect 546162 219922 546218 219978
rect 561250 220294 561306 220350
rect 561374 220294 561430 220350
rect 561498 220294 561554 220350
rect 561622 220294 561678 220350
rect 561250 220170 561306 220226
rect 561374 220170 561430 220226
rect 561498 220170 561554 220226
rect 561622 220170 561678 220226
rect 561250 220046 561306 220102
rect 561374 220046 561430 220102
rect 561498 220046 561554 220102
rect 561622 220046 561678 220102
rect 561250 219922 561306 219978
rect 561374 219922 561430 219978
rect 561498 219922 561554 219978
rect 561622 219922 561678 219978
rect 131318 208294 131374 208350
rect 131442 208294 131498 208350
rect 131318 208170 131374 208226
rect 131442 208170 131498 208226
rect 131318 208046 131374 208102
rect 131442 208046 131498 208102
rect 131318 207922 131374 207978
rect 131442 207922 131498 207978
rect 162038 208294 162094 208350
rect 162162 208294 162218 208350
rect 162038 208170 162094 208226
rect 162162 208170 162218 208226
rect 162038 208046 162094 208102
rect 162162 208046 162218 208102
rect 162038 207922 162094 207978
rect 162162 207922 162218 207978
rect 192758 208294 192814 208350
rect 192882 208294 192938 208350
rect 192758 208170 192814 208226
rect 192882 208170 192938 208226
rect 192758 208046 192814 208102
rect 192882 208046 192938 208102
rect 192758 207922 192814 207978
rect 192882 207922 192938 207978
rect 223478 208294 223534 208350
rect 223602 208294 223658 208350
rect 223478 208170 223534 208226
rect 223602 208170 223658 208226
rect 223478 208046 223534 208102
rect 223602 208046 223658 208102
rect 223478 207922 223534 207978
rect 223602 207922 223658 207978
rect 254198 208294 254254 208350
rect 254322 208294 254378 208350
rect 254198 208170 254254 208226
rect 254322 208170 254378 208226
rect 254198 208046 254254 208102
rect 254322 208046 254378 208102
rect 254198 207922 254254 207978
rect 254322 207922 254378 207978
rect 284918 208294 284974 208350
rect 285042 208294 285098 208350
rect 284918 208170 284974 208226
rect 285042 208170 285098 208226
rect 284918 208046 284974 208102
rect 285042 208046 285098 208102
rect 284918 207922 284974 207978
rect 285042 207922 285098 207978
rect 315638 208294 315694 208350
rect 315762 208294 315818 208350
rect 315638 208170 315694 208226
rect 315762 208170 315818 208226
rect 315638 208046 315694 208102
rect 315762 208046 315818 208102
rect 315638 207922 315694 207978
rect 315762 207922 315818 207978
rect 346358 208294 346414 208350
rect 346482 208294 346538 208350
rect 346358 208170 346414 208226
rect 346482 208170 346538 208226
rect 346358 208046 346414 208102
rect 346482 208046 346538 208102
rect 346358 207922 346414 207978
rect 346482 207922 346538 207978
rect 377078 208294 377134 208350
rect 377202 208294 377258 208350
rect 377078 208170 377134 208226
rect 377202 208170 377258 208226
rect 377078 208046 377134 208102
rect 377202 208046 377258 208102
rect 377078 207922 377134 207978
rect 377202 207922 377258 207978
rect 407798 208294 407854 208350
rect 407922 208294 407978 208350
rect 407798 208170 407854 208226
rect 407922 208170 407978 208226
rect 407798 208046 407854 208102
rect 407922 208046 407978 208102
rect 407798 207922 407854 207978
rect 407922 207922 407978 207978
rect 438518 208294 438574 208350
rect 438642 208294 438698 208350
rect 438518 208170 438574 208226
rect 438642 208170 438698 208226
rect 438518 208046 438574 208102
rect 438642 208046 438698 208102
rect 438518 207922 438574 207978
rect 438642 207922 438698 207978
rect 469238 208294 469294 208350
rect 469362 208294 469418 208350
rect 469238 208170 469294 208226
rect 469362 208170 469418 208226
rect 469238 208046 469294 208102
rect 469362 208046 469418 208102
rect 469238 207922 469294 207978
rect 469362 207922 469418 207978
rect 499958 208294 500014 208350
rect 500082 208294 500138 208350
rect 499958 208170 500014 208226
rect 500082 208170 500138 208226
rect 499958 208046 500014 208102
rect 500082 208046 500138 208102
rect 499958 207922 500014 207978
rect 500082 207922 500138 207978
rect 530678 208294 530734 208350
rect 530802 208294 530858 208350
rect 530678 208170 530734 208226
rect 530802 208170 530858 208226
rect 530678 208046 530734 208102
rect 530802 208046 530858 208102
rect 530678 207922 530734 207978
rect 530802 207922 530858 207978
rect 111250 202294 111306 202350
rect 111374 202294 111430 202350
rect 111498 202294 111554 202350
rect 111622 202294 111678 202350
rect 111250 202170 111306 202226
rect 111374 202170 111430 202226
rect 111498 202170 111554 202226
rect 111622 202170 111678 202226
rect 111250 202046 111306 202102
rect 111374 202046 111430 202102
rect 111498 202046 111554 202102
rect 111622 202046 111678 202102
rect 111250 201922 111306 201978
rect 111374 201922 111430 201978
rect 111498 201922 111554 201978
rect 111622 201922 111678 201978
rect 96970 190294 97026 190350
rect 97094 190294 97150 190350
rect 97218 190294 97274 190350
rect 97342 190294 97398 190350
rect 96970 190170 97026 190226
rect 97094 190170 97150 190226
rect 97218 190170 97274 190226
rect 97342 190170 97398 190226
rect 96970 190046 97026 190102
rect 97094 190046 97150 190102
rect 97218 190046 97274 190102
rect 97342 190046 97398 190102
rect 96970 189922 97026 189978
rect 97094 189922 97150 189978
rect 97218 189922 97274 189978
rect 97342 189922 97398 189978
rect 100598 190294 100654 190350
rect 100722 190294 100778 190350
rect 100598 190170 100654 190226
rect 100722 190170 100778 190226
rect 100598 190046 100654 190102
rect 100722 190046 100778 190102
rect 100598 189922 100654 189978
rect 100722 189922 100778 189978
rect 115958 202294 116014 202350
rect 116082 202294 116138 202350
rect 115958 202170 116014 202226
rect 116082 202170 116138 202226
rect 115958 202046 116014 202102
rect 116082 202046 116138 202102
rect 115958 201922 116014 201978
rect 116082 201922 116138 201978
rect 146678 202294 146734 202350
rect 146802 202294 146858 202350
rect 146678 202170 146734 202226
rect 146802 202170 146858 202226
rect 146678 202046 146734 202102
rect 146802 202046 146858 202102
rect 146678 201922 146734 201978
rect 146802 201922 146858 201978
rect 177398 202294 177454 202350
rect 177522 202294 177578 202350
rect 177398 202170 177454 202226
rect 177522 202170 177578 202226
rect 177398 202046 177454 202102
rect 177522 202046 177578 202102
rect 177398 201922 177454 201978
rect 177522 201922 177578 201978
rect 208118 202294 208174 202350
rect 208242 202294 208298 202350
rect 208118 202170 208174 202226
rect 208242 202170 208298 202226
rect 208118 202046 208174 202102
rect 208242 202046 208298 202102
rect 208118 201922 208174 201978
rect 208242 201922 208298 201978
rect 238838 202294 238894 202350
rect 238962 202294 239018 202350
rect 238838 202170 238894 202226
rect 238962 202170 239018 202226
rect 238838 202046 238894 202102
rect 238962 202046 239018 202102
rect 238838 201922 238894 201978
rect 238962 201922 239018 201978
rect 269558 202294 269614 202350
rect 269682 202294 269738 202350
rect 269558 202170 269614 202226
rect 269682 202170 269738 202226
rect 269558 202046 269614 202102
rect 269682 202046 269738 202102
rect 269558 201922 269614 201978
rect 269682 201922 269738 201978
rect 300278 202294 300334 202350
rect 300402 202294 300458 202350
rect 300278 202170 300334 202226
rect 300402 202170 300458 202226
rect 300278 202046 300334 202102
rect 300402 202046 300458 202102
rect 300278 201922 300334 201978
rect 300402 201922 300458 201978
rect 330998 202294 331054 202350
rect 331122 202294 331178 202350
rect 330998 202170 331054 202226
rect 331122 202170 331178 202226
rect 330998 202046 331054 202102
rect 331122 202046 331178 202102
rect 330998 201922 331054 201978
rect 331122 201922 331178 201978
rect 361718 202294 361774 202350
rect 361842 202294 361898 202350
rect 361718 202170 361774 202226
rect 361842 202170 361898 202226
rect 361718 202046 361774 202102
rect 361842 202046 361898 202102
rect 361718 201922 361774 201978
rect 361842 201922 361898 201978
rect 392438 202294 392494 202350
rect 392562 202294 392618 202350
rect 392438 202170 392494 202226
rect 392562 202170 392618 202226
rect 392438 202046 392494 202102
rect 392562 202046 392618 202102
rect 392438 201922 392494 201978
rect 392562 201922 392618 201978
rect 423158 202294 423214 202350
rect 423282 202294 423338 202350
rect 423158 202170 423214 202226
rect 423282 202170 423338 202226
rect 423158 202046 423214 202102
rect 423282 202046 423338 202102
rect 423158 201922 423214 201978
rect 423282 201922 423338 201978
rect 453878 202294 453934 202350
rect 454002 202294 454058 202350
rect 453878 202170 453934 202226
rect 454002 202170 454058 202226
rect 453878 202046 453934 202102
rect 454002 202046 454058 202102
rect 453878 201922 453934 201978
rect 454002 201922 454058 201978
rect 484598 202294 484654 202350
rect 484722 202294 484778 202350
rect 484598 202170 484654 202226
rect 484722 202170 484778 202226
rect 484598 202046 484654 202102
rect 484722 202046 484778 202102
rect 484598 201922 484654 201978
rect 484722 201922 484778 201978
rect 515318 202294 515374 202350
rect 515442 202294 515498 202350
rect 515318 202170 515374 202226
rect 515442 202170 515498 202226
rect 515318 202046 515374 202102
rect 515442 202046 515498 202102
rect 515318 201922 515374 201978
rect 515442 201922 515498 201978
rect 546038 202294 546094 202350
rect 546162 202294 546218 202350
rect 546038 202170 546094 202226
rect 546162 202170 546218 202226
rect 546038 202046 546094 202102
rect 546162 202046 546218 202102
rect 546038 201922 546094 201978
rect 546162 201922 546218 201978
rect 561250 202294 561306 202350
rect 561374 202294 561430 202350
rect 561498 202294 561554 202350
rect 561622 202294 561678 202350
rect 561250 202170 561306 202226
rect 561374 202170 561430 202226
rect 561498 202170 561554 202226
rect 561622 202170 561678 202226
rect 561250 202046 561306 202102
rect 561374 202046 561430 202102
rect 561498 202046 561554 202102
rect 561622 202046 561678 202102
rect 561250 201922 561306 201978
rect 561374 201922 561430 201978
rect 561498 201922 561554 201978
rect 561622 201922 561678 201978
rect 131318 190294 131374 190350
rect 131442 190294 131498 190350
rect 131318 190170 131374 190226
rect 131442 190170 131498 190226
rect 131318 190046 131374 190102
rect 131442 190046 131498 190102
rect 131318 189922 131374 189978
rect 131442 189922 131498 189978
rect 162038 190294 162094 190350
rect 162162 190294 162218 190350
rect 162038 190170 162094 190226
rect 162162 190170 162218 190226
rect 162038 190046 162094 190102
rect 162162 190046 162218 190102
rect 162038 189922 162094 189978
rect 162162 189922 162218 189978
rect 192758 190294 192814 190350
rect 192882 190294 192938 190350
rect 192758 190170 192814 190226
rect 192882 190170 192938 190226
rect 192758 190046 192814 190102
rect 192882 190046 192938 190102
rect 192758 189922 192814 189978
rect 192882 189922 192938 189978
rect 223478 190294 223534 190350
rect 223602 190294 223658 190350
rect 223478 190170 223534 190226
rect 223602 190170 223658 190226
rect 223478 190046 223534 190102
rect 223602 190046 223658 190102
rect 223478 189922 223534 189978
rect 223602 189922 223658 189978
rect 254198 190294 254254 190350
rect 254322 190294 254378 190350
rect 254198 190170 254254 190226
rect 254322 190170 254378 190226
rect 254198 190046 254254 190102
rect 254322 190046 254378 190102
rect 254198 189922 254254 189978
rect 254322 189922 254378 189978
rect 284918 190294 284974 190350
rect 285042 190294 285098 190350
rect 284918 190170 284974 190226
rect 285042 190170 285098 190226
rect 284918 190046 284974 190102
rect 285042 190046 285098 190102
rect 284918 189922 284974 189978
rect 285042 189922 285098 189978
rect 315638 190294 315694 190350
rect 315762 190294 315818 190350
rect 315638 190170 315694 190226
rect 315762 190170 315818 190226
rect 315638 190046 315694 190102
rect 315762 190046 315818 190102
rect 315638 189922 315694 189978
rect 315762 189922 315818 189978
rect 346358 190294 346414 190350
rect 346482 190294 346538 190350
rect 346358 190170 346414 190226
rect 346482 190170 346538 190226
rect 346358 190046 346414 190102
rect 346482 190046 346538 190102
rect 346358 189922 346414 189978
rect 346482 189922 346538 189978
rect 377078 190294 377134 190350
rect 377202 190294 377258 190350
rect 377078 190170 377134 190226
rect 377202 190170 377258 190226
rect 377078 190046 377134 190102
rect 377202 190046 377258 190102
rect 377078 189922 377134 189978
rect 377202 189922 377258 189978
rect 407798 190294 407854 190350
rect 407922 190294 407978 190350
rect 407798 190170 407854 190226
rect 407922 190170 407978 190226
rect 407798 190046 407854 190102
rect 407922 190046 407978 190102
rect 407798 189922 407854 189978
rect 407922 189922 407978 189978
rect 438518 190294 438574 190350
rect 438642 190294 438698 190350
rect 438518 190170 438574 190226
rect 438642 190170 438698 190226
rect 438518 190046 438574 190102
rect 438642 190046 438698 190102
rect 438518 189922 438574 189978
rect 438642 189922 438698 189978
rect 469238 190294 469294 190350
rect 469362 190294 469418 190350
rect 469238 190170 469294 190226
rect 469362 190170 469418 190226
rect 469238 190046 469294 190102
rect 469362 190046 469418 190102
rect 469238 189922 469294 189978
rect 469362 189922 469418 189978
rect 499958 190294 500014 190350
rect 500082 190294 500138 190350
rect 499958 190170 500014 190226
rect 500082 190170 500138 190226
rect 499958 190046 500014 190102
rect 500082 190046 500138 190102
rect 499958 189922 500014 189978
rect 500082 189922 500138 189978
rect 530678 190294 530734 190350
rect 530802 190294 530858 190350
rect 530678 190170 530734 190226
rect 530802 190170 530858 190226
rect 530678 190046 530734 190102
rect 530802 190046 530858 190102
rect 530678 189922 530734 189978
rect 530802 189922 530858 189978
rect 111250 184294 111306 184350
rect 111374 184294 111430 184350
rect 111498 184294 111554 184350
rect 111622 184294 111678 184350
rect 111250 184170 111306 184226
rect 111374 184170 111430 184226
rect 111498 184170 111554 184226
rect 111622 184170 111678 184226
rect 111250 184046 111306 184102
rect 111374 184046 111430 184102
rect 111498 184046 111554 184102
rect 111622 184046 111678 184102
rect 111250 183922 111306 183978
rect 111374 183922 111430 183978
rect 111498 183922 111554 183978
rect 111622 183922 111678 183978
rect 96970 172294 97026 172350
rect 97094 172294 97150 172350
rect 97218 172294 97274 172350
rect 97342 172294 97398 172350
rect 96970 172170 97026 172226
rect 97094 172170 97150 172226
rect 97218 172170 97274 172226
rect 97342 172170 97398 172226
rect 96970 172046 97026 172102
rect 97094 172046 97150 172102
rect 97218 172046 97274 172102
rect 97342 172046 97398 172102
rect 96970 171922 97026 171978
rect 97094 171922 97150 171978
rect 97218 171922 97274 171978
rect 97342 171922 97398 171978
rect 100598 172294 100654 172350
rect 100722 172294 100778 172350
rect 100598 172170 100654 172226
rect 100722 172170 100778 172226
rect 100598 172046 100654 172102
rect 100722 172046 100778 172102
rect 100598 171922 100654 171978
rect 100722 171922 100778 171978
rect 115958 184294 116014 184350
rect 116082 184294 116138 184350
rect 115958 184170 116014 184226
rect 116082 184170 116138 184226
rect 115958 184046 116014 184102
rect 116082 184046 116138 184102
rect 115958 183922 116014 183978
rect 116082 183922 116138 183978
rect 146678 184294 146734 184350
rect 146802 184294 146858 184350
rect 146678 184170 146734 184226
rect 146802 184170 146858 184226
rect 146678 184046 146734 184102
rect 146802 184046 146858 184102
rect 146678 183922 146734 183978
rect 146802 183922 146858 183978
rect 177398 184294 177454 184350
rect 177522 184294 177578 184350
rect 177398 184170 177454 184226
rect 177522 184170 177578 184226
rect 177398 184046 177454 184102
rect 177522 184046 177578 184102
rect 177398 183922 177454 183978
rect 177522 183922 177578 183978
rect 208118 184294 208174 184350
rect 208242 184294 208298 184350
rect 208118 184170 208174 184226
rect 208242 184170 208298 184226
rect 208118 184046 208174 184102
rect 208242 184046 208298 184102
rect 208118 183922 208174 183978
rect 208242 183922 208298 183978
rect 238838 184294 238894 184350
rect 238962 184294 239018 184350
rect 238838 184170 238894 184226
rect 238962 184170 239018 184226
rect 238838 184046 238894 184102
rect 238962 184046 239018 184102
rect 238838 183922 238894 183978
rect 238962 183922 239018 183978
rect 269558 184294 269614 184350
rect 269682 184294 269738 184350
rect 269558 184170 269614 184226
rect 269682 184170 269738 184226
rect 269558 184046 269614 184102
rect 269682 184046 269738 184102
rect 269558 183922 269614 183978
rect 269682 183922 269738 183978
rect 300278 184294 300334 184350
rect 300402 184294 300458 184350
rect 300278 184170 300334 184226
rect 300402 184170 300458 184226
rect 300278 184046 300334 184102
rect 300402 184046 300458 184102
rect 300278 183922 300334 183978
rect 300402 183922 300458 183978
rect 330998 184294 331054 184350
rect 331122 184294 331178 184350
rect 330998 184170 331054 184226
rect 331122 184170 331178 184226
rect 330998 184046 331054 184102
rect 331122 184046 331178 184102
rect 330998 183922 331054 183978
rect 331122 183922 331178 183978
rect 361718 184294 361774 184350
rect 361842 184294 361898 184350
rect 361718 184170 361774 184226
rect 361842 184170 361898 184226
rect 361718 184046 361774 184102
rect 361842 184046 361898 184102
rect 361718 183922 361774 183978
rect 361842 183922 361898 183978
rect 392438 184294 392494 184350
rect 392562 184294 392618 184350
rect 392438 184170 392494 184226
rect 392562 184170 392618 184226
rect 392438 184046 392494 184102
rect 392562 184046 392618 184102
rect 392438 183922 392494 183978
rect 392562 183922 392618 183978
rect 423158 184294 423214 184350
rect 423282 184294 423338 184350
rect 423158 184170 423214 184226
rect 423282 184170 423338 184226
rect 423158 184046 423214 184102
rect 423282 184046 423338 184102
rect 423158 183922 423214 183978
rect 423282 183922 423338 183978
rect 453878 184294 453934 184350
rect 454002 184294 454058 184350
rect 453878 184170 453934 184226
rect 454002 184170 454058 184226
rect 453878 184046 453934 184102
rect 454002 184046 454058 184102
rect 453878 183922 453934 183978
rect 454002 183922 454058 183978
rect 484598 184294 484654 184350
rect 484722 184294 484778 184350
rect 484598 184170 484654 184226
rect 484722 184170 484778 184226
rect 484598 184046 484654 184102
rect 484722 184046 484778 184102
rect 484598 183922 484654 183978
rect 484722 183922 484778 183978
rect 515318 184294 515374 184350
rect 515442 184294 515498 184350
rect 515318 184170 515374 184226
rect 515442 184170 515498 184226
rect 515318 184046 515374 184102
rect 515442 184046 515498 184102
rect 515318 183922 515374 183978
rect 515442 183922 515498 183978
rect 546038 184294 546094 184350
rect 546162 184294 546218 184350
rect 546038 184170 546094 184226
rect 546162 184170 546218 184226
rect 546038 184046 546094 184102
rect 546162 184046 546218 184102
rect 546038 183922 546094 183978
rect 546162 183922 546218 183978
rect 561250 184294 561306 184350
rect 561374 184294 561430 184350
rect 561498 184294 561554 184350
rect 561622 184294 561678 184350
rect 561250 184170 561306 184226
rect 561374 184170 561430 184226
rect 561498 184170 561554 184226
rect 561622 184170 561678 184226
rect 561250 184046 561306 184102
rect 561374 184046 561430 184102
rect 561498 184046 561554 184102
rect 561622 184046 561678 184102
rect 561250 183922 561306 183978
rect 561374 183922 561430 183978
rect 561498 183922 561554 183978
rect 561622 183922 561678 183978
rect 131318 172294 131374 172350
rect 131442 172294 131498 172350
rect 131318 172170 131374 172226
rect 131442 172170 131498 172226
rect 131318 172046 131374 172102
rect 131442 172046 131498 172102
rect 131318 171922 131374 171978
rect 131442 171922 131498 171978
rect 162038 172294 162094 172350
rect 162162 172294 162218 172350
rect 162038 172170 162094 172226
rect 162162 172170 162218 172226
rect 162038 172046 162094 172102
rect 162162 172046 162218 172102
rect 162038 171922 162094 171978
rect 162162 171922 162218 171978
rect 192758 172294 192814 172350
rect 192882 172294 192938 172350
rect 192758 172170 192814 172226
rect 192882 172170 192938 172226
rect 192758 172046 192814 172102
rect 192882 172046 192938 172102
rect 192758 171922 192814 171978
rect 192882 171922 192938 171978
rect 223478 172294 223534 172350
rect 223602 172294 223658 172350
rect 223478 172170 223534 172226
rect 223602 172170 223658 172226
rect 223478 172046 223534 172102
rect 223602 172046 223658 172102
rect 223478 171922 223534 171978
rect 223602 171922 223658 171978
rect 254198 172294 254254 172350
rect 254322 172294 254378 172350
rect 254198 172170 254254 172226
rect 254322 172170 254378 172226
rect 254198 172046 254254 172102
rect 254322 172046 254378 172102
rect 254198 171922 254254 171978
rect 254322 171922 254378 171978
rect 284918 172294 284974 172350
rect 285042 172294 285098 172350
rect 284918 172170 284974 172226
rect 285042 172170 285098 172226
rect 284918 172046 284974 172102
rect 285042 172046 285098 172102
rect 284918 171922 284974 171978
rect 285042 171922 285098 171978
rect 315638 172294 315694 172350
rect 315762 172294 315818 172350
rect 315638 172170 315694 172226
rect 315762 172170 315818 172226
rect 315638 172046 315694 172102
rect 315762 172046 315818 172102
rect 315638 171922 315694 171978
rect 315762 171922 315818 171978
rect 346358 172294 346414 172350
rect 346482 172294 346538 172350
rect 346358 172170 346414 172226
rect 346482 172170 346538 172226
rect 346358 172046 346414 172102
rect 346482 172046 346538 172102
rect 346358 171922 346414 171978
rect 346482 171922 346538 171978
rect 377078 172294 377134 172350
rect 377202 172294 377258 172350
rect 377078 172170 377134 172226
rect 377202 172170 377258 172226
rect 377078 172046 377134 172102
rect 377202 172046 377258 172102
rect 377078 171922 377134 171978
rect 377202 171922 377258 171978
rect 407798 172294 407854 172350
rect 407922 172294 407978 172350
rect 407798 172170 407854 172226
rect 407922 172170 407978 172226
rect 407798 172046 407854 172102
rect 407922 172046 407978 172102
rect 407798 171922 407854 171978
rect 407922 171922 407978 171978
rect 438518 172294 438574 172350
rect 438642 172294 438698 172350
rect 438518 172170 438574 172226
rect 438642 172170 438698 172226
rect 438518 172046 438574 172102
rect 438642 172046 438698 172102
rect 438518 171922 438574 171978
rect 438642 171922 438698 171978
rect 469238 172294 469294 172350
rect 469362 172294 469418 172350
rect 469238 172170 469294 172226
rect 469362 172170 469418 172226
rect 469238 172046 469294 172102
rect 469362 172046 469418 172102
rect 469238 171922 469294 171978
rect 469362 171922 469418 171978
rect 499958 172294 500014 172350
rect 500082 172294 500138 172350
rect 499958 172170 500014 172226
rect 500082 172170 500138 172226
rect 499958 172046 500014 172102
rect 500082 172046 500138 172102
rect 499958 171922 500014 171978
rect 500082 171922 500138 171978
rect 530678 172294 530734 172350
rect 530802 172294 530858 172350
rect 530678 172170 530734 172226
rect 530802 172170 530858 172226
rect 530678 172046 530734 172102
rect 530802 172046 530858 172102
rect 530678 171922 530734 171978
rect 530802 171922 530858 171978
rect 111250 166294 111306 166350
rect 111374 166294 111430 166350
rect 111498 166294 111554 166350
rect 111622 166294 111678 166350
rect 111250 166170 111306 166226
rect 111374 166170 111430 166226
rect 111498 166170 111554 166226
rect 111622 166170 111678 166226
rect 111250 166046 111306 166102
rect 111374 166046 111430 166102
rect 111498 166046 111554 166102
rect 111622 166046 111678 166102
rect 111250 165922 111306 165978
rect 111374 165922 111430 165978
rect 111498 165922 111554 165978
rect 111622 165922 111678 165978
rect 96970 154294 97026 154350
rect 97094 154294 97150 154350
rect 97218 154294 97274 154350
rect 97342 154294 97398 154350
rect 96970 154170 97026 154226
rect 97094 154170 97150 154226
rect 97218 154170 97274 154226
rect 97342 154170 97398 154226
rect 96970 154046 97026 154102
rect 97094 154046 97150 154102
rect 97218 154046 97274 154102
rect 97342 154046 97398 154102
rect 96970 153922 97026 153978
rect 97094 153922 97150 153978
rect 97218 153922 97274 153978
rect 97342 153922 97398 153978
rect 100598 154294 100654 154350
rect 100722 154294 100778 154350
rect 100598 154170 100654 154226
rect 100722 154170 100778 154226
rect 100598 154046 100654 154102
rect 100722 154046 100778 154102
rect 100598 153922 100654 153978
rect 100722 153922 100778 153978
rect 115958 166294 116014 166350
rect 116082 166294 116138 166350
rect 115958 166170 116014 166226
rect 116082 166170 116138 166226
rect 115958 166046 116014 166102
rect 116082 166046 116138 166102
rect 115958 165922 116014 165978
rect 116082 165922 116138 165978
rect 146678 166294 146734 166350
rect 146802 166294 146858 166350
rect 146678 166170 146734 166226
rect 146802 166170 146858 166226
rect 146678 166046 146734 166102
rect 146802 166046 146858 166102
rect 146678 165922 146734 165978
rect 146802 165922 146858 165978
rect 177398 166294 177454 166350
rect 177522 166294 177578 166350
rect 177398 166170 177454 166226
rect 177522 166170 177578 166226
rect 177398 166046 177454 166102
rect 177522 166046 177578 166102
rect 177398 165922 177454 165978
rect 177522 165922 177578 165978
rect 208118 166294 208174 166350
rect 208242 166294 208298 166350
rect 208118 166170 208174 166226
rect 208242 166170 208298 166226
rect 208118 166046 208174 166102
rect 208242 166046 208298 166102
rect 208118 165922 208174 165978
rect 208242 165922 208298 165978
rect 238838 166294 238894 166350
rect 238962 166294 239018 166350
rect 238838 166170 238894 166226
rect 238962 166170 239018 166226
rect 238838 166046 238894 166102
rect 238962 166046 239018 166102
rect 238838 165922 238894 165978
rect 238962 165922 239018 165978
rect 269558 166294 269614 166350
rect 269682 166294 269738 166350
rect 269558 166170 269614 166226
rect 269682 166170 269738 166226
rect 269558 166046 269614 166102
rect 269682 166046 269738 166102
rect 269558 165922 269614 165978
rect 269682 165922 269738 165978
rect 300278 166294 300334 166350
rect 300402 166294 300458 166350
rect 300278 166170 300334 166226
rect 300402 166170 300458 166226
rect 300278 166046 300334 166102
rect 300402 166046 300458 166102
rect 300278 165922 300334 165978
rect 300402 165922 300458 165978
rect 330998 166294 331054 166350
rect 331122 166294 331178 166350
rect 330998 166170 331054 166226
rect 331122 166170 331178 166226
rect 330998 166046 331054 166102
rect 331122 166046 331178 166102
rect 330998 165922 331054 165978
rect 331122 165922 331178 165978
rect 361718 166294 361774 166350
rect 361842 166294 361898 166350
rect 361718 166170 361774 166226
rect 361842 166170 361898 166226
rect 361718 166046 361774 166102
rect 361842 166046 361898 166102
rect 361718 165922 361774 165978
rect 361842 165922 361898 165978
rect 392438 166294 392494 166350
rect 392562 166294 392618 166350
rect 392438 166170 392494 166226
rect 392562 166170 392618 166226
rect 392438 166046 392494 166102
rect 392562 166046 392618 166102
rect 392438 165922 392494 165978
rect 392562 165922 392618 165978
rect 423158 166294 423214 166350
rect 423282 166294 423338 166350
rect 423158 166170 423214 166226
rect 423282 166170 423338 166226
rect 423158 166046 423214 166102
rect 423282 166046 423338 166102
rect 423158 165922 423214 165978
rect 423282 165922 423338 165978
rect 453878 166294 453934 166350
rect 454002 166294 454058 166350
rect 453878 166170 453934 166226
rect 454002 166170 454058 166226
rect 453878 166046 453934 166102
rect 454002 166046 454058 166102
rect 453878 165922 453934 165978
rect 454002 165922 454058 165978
rect 484598 166294 484654 166350
rect 484722 166294 484778 166350
rect 484598 166170 484654 166226
rect 484722 166170 484778 166226
rect 484598 166046 484654 166102
rect 484722 166046 484778 166102
rect 484598 165922 484654 165978
rect 484722 165922 484778 165978
rect 515318 166294 515374 166350
rect 515442 166294 515498 166350
rect 515318 166170 515374 166226
rect 515442 166170 515498 166226
rect 515318 166046 515374 166102
rect 515442 166046 515498 166102
rect 515318 165922 515374 165978
rect 515442 165922 515498 165978
rect 546038 166294 546094 166350
rect 546162 166294 546218 166350
rect 546038 166170 546094 166226
rect 546162 166170 546218 166226
rect 546038 166046 546094 166102
rect 546162 166046 546218 166102
rect 546038 165922 546094 165978
rect 546162 165922 546218 165978
rect 561250 166294 561306 166350
rect 561374 166294 561430 166350
rect 561498 166294 561554 166350
rect 561622 166294 561678 166350
rect 561250 166170 561306 166226
rect 561374 166170 561430 166226
rect 561498 166170 561554 166226
rect 561622 166170 561678 166226
rect 561250 166046 561306 166102
rect 561374 166046 561430 166102
rect 561498 166046 561554 166102
rect 561622 166046 561678 166102
rect 561250 165922 561306 165978
rect 561374 165922 561430 165978
rect 561498 165922 561554 165978
rect 561622 165922 561678 165978
rect 131318 154294 131374 154350
rect 131442 154294 131498 154350
rect 131318 154170 131374 154226
rect 131442 154170 131498 154226
rect 131318 154046 131374 154102
rect 131442 154046 131498 154102
rect 131318 153922 131374 153978
rect 131442 153922 131498 153978
rect 162038 154294 162094 154350
rect 162162 154294 162218 154350
rect 162038 154170 162094 154226
rect 162162 154170 162218 154226
rect 162038 154046 162094 154102
rect 162162 154046 162218 154102
rect 162038 153922 162094 153978
rect 162162 153922 162218 153978
rect 192758 154294 192814 154350
rect 192882 154294 192938 154350
rect 192758 154170 192814 154226
rect 192882 154170 192938 154226
rect 192758 154046 192814 154102
rect 192882 154046 192938 154102
rect 192758 153922 192814 153978
rect 192882 153922 192938 153978
rect 223478 154294 223534 154350
rect 223602 154294 223658 154350
rect 223478 154170 223534 154226
rect 223602 154170 223658 154226
rect 223478 154046 223534 154102
rect 223602 154046 223658 154102
rect 223478 153922 223534 153978
rect 223602 153922 223658 153978
rect 254198 154294 254254 154350
rect 254322 154294 254378 154350
rect 254198 154170 254254 154226
rect 254322 154170 254378 154226
rect 254198 154046 254254 154102
rect 254322 154046 254378 154102
rect 254198 153922 254254 153978
rect 254322 153922 254378 153978
rect 284918 154294 284974 154350
rect 285042 154294 285098 154350
rect 284918 154170 284974 154226
rect 285042 154170 285098 154226
rect 284918 154046 284974 154102
rect 285042 154046 285098 154102
rect 284918 153922 284974 153978
rect 285042 153922 285098 153978
rect 315638 154294 315694 154350
rect 315762 154294 315818 154350
rect 315638 154170 315694 154226
rect 315762 154170 315818 154226
rect 315638 154046 315694 154102
rect 315762 154046 315818 154102
rect 315638 153922 315694 153978
rect 315762 153922 315818 153978
rect 346358 154294 346414 154350
rect 346482 154294 346538 154350
rect 346358 154170 346414 154226
rect 346482 154170 346538 154226
rect 346358 154046 346414 154102
rect 346482 154046 346538 154102
rect 346358 153922 346414 153978
rect 346482 153922 346538 153978
rect 377078 154294 377134 154350
rect 377202 154294 377258 154350
rect 377078 154170 377134 154226
rect 377202 154170 377258 154226
rect 377078 154046 377134 154102
rect 377202 154046 377258 154102
rect 377078 153922 377134 153978
rect 377202 153922 377258 153978
rect 407798 154294 407854 154350
rect 407922 154294 407978 154350
rect 407798 154170 407854 154226
rect 407922 154170 407978 154226
rect 407798 154046 407854 154102
rect 407922 154046 407978 154102
rect 407798 153922 407854 153978
rect 407922 153922 407978 153978
rect 438518 154294 438574 154350
rect 438642 154294 438698 154350
rect 438518 154170 438574 154226
rect 438642 154170 438698 154226
rect 438518 154046 438574 154102
rect 438642 154046 438698 154102
rect 438518 153922 438574 153978
rect 438642 153922 438698 153978
rect 469238 154294 469294 154350
rect 469362 154294 469418 154350
rect 469238 154170 469294 154226
rect 469362 154170 469418 154226
rect 469238 154046 469294 154102
rect 469362 154046 469418 154102
rect 469238 153922 469294 153978
rect 469362 153922 469418 153978
rect 499958 154294 500014 154350
rect 500082 154294 500138 154350
rect 499958 154170 500014 154226
rect 500082 154170 500138 154226
rect 499958 154046 500014 154102
rect 500082 154046 500138 154102
rect 499958 153922 500014 153978
rect 500082 153922 500138 153978
rect 530678 154294 530734 154350
rect 530802 154294 530858 154350
rect 530678 154170 530734 154226
rect 530802 154170 530858 154226
rect 530678 154046 530734 154102
rect 530802 154046 530858 154102
rect 530678 153922 530734 153978
rect 530802 153922 530858 153978
rect 111250 148294 111306 148350
rect 111374 148294 111430 148350
rect 111498 148294 111554 148350
rect 111622 148294 111678 148350
rect 111250 148170 111306 148226
rect 111374 148170 111430 148226
rect 111498 148170 111554 148226
rect 111622 148170 111678 148226
rect 111250 148046 111306 148102
rect 111374 148046 111430 148102
rect 111498 148046 111554 148102
rect 111622 148046 111678 148102
rect 111250 147922 111306 147978
rect 111374 147922 111430 147978
rect 111498 147922 111554 147978
rect 111622 147922 111678 147978
rect 96970 136294 97026 136350
rect 97094 136294 97150 136350
rect 97218 136294 97274 136350
rect 97342 136294 97398 136350
rect 96970 136170 97026 136226
rect 97094 136170 97150 136226
rect 97218 136170 97274 136226
rect 97342 136170 97398 136226
rect 96970 136046 97026 136102
rect 97094 136046 97150 136102
rect 97218 136046 97274 136102
rect 97342 136046 97398 136102
rect 96970 135922 97026 135978
rect 97094 135922 97150 135978
rect 97218 135922 97274 135978
rect 97342 135922 97398 135978
rect 100598 136294 100654 136350
rect 100722 136294 100778 136350
rect 100598 136170 100654 136226
rect 100722 136170 100778 136226
rect 100598 136046 100654 136102
rect 100722 136046 100778 136102
rect 100598 135922 100654 135978
rect 100722 135922 100778 135978
rect 115958 148294 116014 148350
rect 116082 148294 116138 148350
rect 115958 148170 116014 148226
rect 116082 148170 116138 148226
rect 115958 148046 116014 148102
rect 116082 148046 116138 148102
rect 115958 147922 116014 147978
rect 116082 147922 116138 147978
rect 146678 148294 146734 148350
rect 146802 148294 146858 148350
rect 146678 148170 146734 148226
rect 146802 148170 146858 148226
rect 146678 148046 146734 148102
rect 146802 148046 146858 148102
rect 146678 147922 146734 147978
rect 146802 147922 146858 147978
rect 177398 148294 177454 148350
rect 177522 148294 177578 148350
rect 177398 148170 177454 148226
rect 177522 148170 177578 148226
rect 177398 148046 177454 148102
rect 177522 148046 177578 148102
rect 177398 147922 177454 147978
rect 177522 147922 177578 147978
rect 208118 148294 208174 148350
rect 208242 148294 208298 148350
rect 208118 148170 208174 148226
rect 208242 148170 208298 148226
rect 208118 148046 208174 148102
rect 208242 148046 208298 148102
rect 208118 147922 208174 147978
rect 208242 147922 208298 147978
rect 238838 148294 238894 148350
rect 238962 148294 239018 148350
rect 238838 148170 238894 148226
rect 238962 148170 239018 148226
rect 238838 148046 238894 148102
rect 238962 148046 239018 148102
rect 238838 147922 238894 147978
rect 238962 147922 239018 147978
rect 269558 148294 269614 148350
rect 269682 148294 269738 148350
rect 269558 148170 269614 148226
rect 269682 148170 269738 148226
rect 269558 148046 269614 148102
rect 269682 148046 269738 148102
rect 269558 147922 269614 147978
rect 269682 147922 269738 147978
rect 300278 148294 300334 148350
rect 300402 148294 300458 148350
rect 300278 148170 300334 148226
rect 300402 148170 300458 148226
rect 300278 148046 300334 148102
rect 300402 148046 300458 148102
rect 300278 147922 300334 147978
rect 300402 147922 300458 147978
rect 330998 148294 331054 148350
rect 331122 148294 331178 148350
rect 330998 148170 331054 148226
rect 331122 148170 331178 148226
rect 330998 148046 331054 148102
rect 331122 148046 331178 148102
rect 330998 147922 331054 147978
rect 331122 147922 331178 147978
rect 361718 148294 361774 148350
rect 361842 148294 361898 148350
rect 361718 148170 361774 148226
rect 361842 148170 361898 148226
rect 361718 148046 361774 148102
rect 361842 148046 361898 148102
rect 361718 147922 361774 147978
rect 361842 147922 361898 147978
rect 392438 148294 392494 148350
rect 392562 148294 392618 148350
rect 392438 148170 392494 148226
rect 392562 148170 392618 148226
rect 392438 148046 392494 148102
rect 392562 148046 392618 148102
rect 392438 147922 392494 147978
rect 392562 147922 392618 147978
rect 423158 148294 423214 148350
rect 423282 148294 423338 148350
rect 423158 148170 423214 148226
rect 423282 148170 423338 148226
rect 423158 148046 423214 148102
rect 423282 148046 423338 148102
rect 423158 147922 423214 147978
rect 423282 147922 423338 147978
rect 453878 148294 453934 148350
rect 454002 148294 454058 148350
rect 453878 148170 453934 148226
rect 454002 148170 454058 148226
rect 453878 148046 453934 148102
rect 454002 148046 454058 148102
rect 453878 147922 453934 147978
rect 454002 147922 454058 147978
rect 484598 148294 484654 148350
rect 484722 148294 484778 148350
rect 484598 148170 484654 148226
rect 484722 148170 484778 148226
rect 484598 148046 484654 148102
rect 484722 148046 484778 148102
rect 484598 147922 484654 147978
rect 484722 147922 484778 147978
rect 515318 148294 515374 148350
rect 515442 148294 515498 148350
rect 515318 148170 515374 148226
rect 515442 148170 515498 148226
rect 515318 148046 515374 148102
rect 515442 148046 515498 148102
rect 515318 147922 515374 147978
rect 515442 147922 515498 147978
rect 546038 148294 546094 148350
rect 546162 148294 546218 148350
rect 546038 148170 546094 148226
rect 546162 148170 546218 148226
rect 546038 148046 546094 148102
rect 546162 148046 546218 148102
rect 546038 147922 546094 147978
rect 546162 147922 546218 147978
rect 561250 148294 561306 148350
rect 561374 148294 561430 148350
rect 561498 148294 561554 148350
rect 561622 148294 561678 148350
rect 561250 148170 561306 148226
rect 561374 148170 561430 148226
rect 561498 148170 561554 148226
rect 561622 148170 561678 148226
rect 561250 148046 561306 148102
rect 561374 148046 561430 148102
rect 561498 148046 561554 148102
rect 561622 148046 561678 148102
rect 561250 147922 561306 147978
rect 561374 147922 561430 147978
rect 561498 147922 561554 147978
rect 561622 147922 561678 147978
rect 131318 136294 131374 136350
rect 131442 136294 131498 136350
rect 131318 136170 131374 136226
rect 131442 136170 131498 136226
rect 131318 136046 131374 136102
rect 131442 136046 131498 136102
rect 131318 135922 131374 135978
rect 131442 135922 131498 135978
rect 162038 136294 162094 136350
rect 162162 136294 162218 136350
rect 162038 136170 162094 136226
rect 162162 136170 162218 136226
rect 162038 136046 162094 136102
rect 162162 136046 162218 136102
rect 162038 135922 162094 135978
rect 162162 135922 162218 135978
rect 192758 136294 192814 136350
rect 192882 136294 192938 136350
rect 192758 136170 192814 136226
rect 192882 136170 192938 136226
rect 192758 136046 192814 136102
rect 192882 136046 192938 136102
rect 192758 135922 192814 135978
rect 192882 135922 192938 135978
rect 223478 136294 223534 136350
rect 223602 136294 223658 136350
rect 223478 136170 223534 136226
rect 223602 136170 223658 136226
rect 223478 136046 223534 136102
rect 223602 136046 223658 136102
rect 223478 135922 223534 135978
rect 223602 135922 223658 135978
rect 254198 136294 254254 136350
rect 254322 136294 254378 136350
rect 254198 136170 254254 136226
rect 254322 136170 254378 136226
rect 254198 136046 254254 136102
rect 254322 136046 254378 136102
rect 254198 135922 254254 135978
rect 254322 135922 254378 135978
rect 284918 136294 284974 136350
rect 285042 136294 285098 136350
rect 284918 136170 284974 136226
rect 285042 136170 285098 136226
rect 284918 136046 284974 136102
rect 285042 136046 285098 136102
rect 284918 135922 284974 135978
rect 285042 135922 285098 135978
rect 315638 136294 315694 136350
rect 315762 136294 315818 136350
rect 315638 136170 315694 136226
rect 315762 136170 315818 136226
rect 315638 136046 315694 136102
rect 315762 136046 315818 136102
rect 315638 135922 315694 135978
rect 315762 135922 315818 135978
rect 346358 136294 346414 136350
rect 346482 136294 346538 136350
rect 346358 136170 346414 136226
rect 346482 136170 346538 136226
rect 346358 136046 346414 136102
rect 346482 136046 346538 136102
rect 346358 135922 346414 135978
rect 346482 135922 346538 135978
rect 377078 136294 377134 136350
rect 377202 136294 377258 136350
rect 377078 136170 377134 136226
rect 377202 136170 377258 136226
rect 377078 136046 377134 136102
rect 377202 136046 377258 136102
rect 377078 135922 377134 135978
rect 377202 135922 377258 135978
rect 407798 136294 407854 136350
rect 407922 136294 407978 136350
rect 407798 136170 407854 136226
rect 407922 136170 407978 136226
rect 407798 136046 407854 136102
rect 407922 136046 407978 136102
rect 407798 135922 407854 135978
rect 407922 135922 407978 135978
rect 438518 136294 438574 136350
rect 438642 136294 438698 136350
rect 438518 136170 438574 136226
rect 438642 136170 438698 136226
rect 438518 136046 438574 136102
rect 438642 136046 438698 136102
rect 438518 135922 438574 135978
rect 438642 135922 438698 135978
rect 469238 136294 469294 136350
rect 469362 136294 469418 136350
rect 469238 136170 469294 136226
rect 469362 136170 469418 136226
rect 469238 136046 469294 136102
rect 469362 136046 469418 136102
rect 469238 135922 469294 135978
rect 469362 135922 469418 135978
rect 499958 136294 500014 136350
rect 500082 136294 500138 136350
rect 499958 136170 500014 136226
rect 500082 136170 500138 136226
rect 499958 136046 500014 136102
rect 500082 136046 500138 136102
rect 499958 135922 500014 135978
rect 500082 135922 500138 135978
rect 530678 136294 530734 136350
rect 530802 136294 530858 136350
rect 530678 136170 530734 136226
rect 530802 136170 530858 136226
rect 530678 136046 530734 136102
rect 530802 136046 530858 136102
rect 530678 135922 530734 135978
rect 530802 135922 530858 135978
rect 111250 130294 111306 130350
rect 111374 130294 111430 130350
rect 111498 130294 111554 130350
rect 111622 130294 111678 130350
rect 111250 130170 111306 130226
rect 111374 130170 111430 130226
rect 111498 130170 111554 130226
rect 111622 130170 111678 130226
rect 111250 130046 111306 130102
rect 111374 130046 111430 130102
rect 111498 130046 111554 130102
rect 111622 130046 111678 130102
rect 111250 129922 111306 129978
rect 111374 129922 111430 129978
rect 111498 129922 111554 129978
rect 111622 129922 111678 129978
rect 96970 118294 97026 118350
rect 97094 118294 97150 118350
rect 97218 118294 97274 118350
rect 97342 118294 97398 118350
rect 96970 118170 97026 118226
rect 97094 118170 97150 118226
rect 97218 118170 97274 118226
rect 97342 118170 97398 118226
rect 96970 118046 97026 118102
rect 97094 118046 97150 118102
rect 97218 118046 97274 118102
rect 97342 118046 97398 118102
rect 96970 117922 97026 117978
rect 97094 117922 97150 117978
rect 97218 117922 97274 117978
rect 97342 117922 97398 117978
rect 100598 118294 100654 118350
rect 100722 118294 100778 118350
rect 100598 118170 100654 118226
rect 100722 118170 100778 118226
rect 100598 118046 100654 118102
rect 100722 118046 100778 118102
rect 100598 117922 100654 117978
rect 100722 117922 100778 117978
rect 115958 130294 116014 130350
rect 116082 130294 116138 130350
rect 115958 130170 116014 130226
rect 116082 130170 116138 130226
rect 115958 130046 116014 130102
rect 116082 130046 116138 130102
rect 115958 129922 116014 129978
rect 116082 129922 116138 129978
rect 146678 130294 146734 130350
rect 146802 130294 146858 130350
rect 146678 130170 146734 130226
rect 146802 130170 146858 130226
rect 146678 130046 146734 130102
rect 146802 130046 146858 130102
rect 146678 129922 146734 129978
rect 146802 129922 146858 129978
rect 177398 130294 177454 130350
rect 177522 130294 177578 130350
rect 177398 130170 177454 130226
rect 177522 130170 177578 130226
rect 177398 130046 177454 130102
rect 177522 130046 177578 130102
rect 177398 129922 177454 129978
rect 177522 129922 177578 129978
rect 208118 130294 208174 130350
rect 208242 130294 208298 130350
rect 208118 130170 208174 130226
rect 208242 130170 208298 130226
rect 208118 130046 208174 130102
rect 208242 130046 208298 130102
rect 208118 129922 208174 129978
rect 208242 129922 208298 129978
rect 238838 130294 238894 130350
rect 238962 130294 239018 130350
rect 238838 130170 238894 130226
rect 238962 130170 239018 130226
rect 238838 130046 238894 130102
rect 238962 130046 239018 130102
rect 238838 129922 238894 129978
rect 238962 129922 239018 129978
rect 269558 130294 269614 130350
rect 269682 130294 269738 130350
rect 269558 130170 269614 130226
rect 269682 130170 269738 130226
rect 269558 130046 269614 130102
rect 269682 130046 269738 130102
rect 269558 129922 269614 129978
rect 269682 129922 269738 129978
rect 300278 130294 300334 130350
rect 300402 130294 300458 130350
rect 300278 130170 300334 130226
rect 300402 130170 300458 130226
rect 300278 130046 300334 130102
rect 300402 130046 300458 130102
rect 300278 129922 300334 129978
rect 300402 129922 300458 129978
rect 330998 130294 331054 130350
rect 331122 130294 331178 130350
rect 330998 130170 331054 130226
rect 331122 130170 331178 130226
rect 330998 130046 331054 130102
rect 331122 130046 331178 130102
rect 330998 129922 331054 129978
rect 331122 129922 331178 129978
rect 361718 130294 361774 130350
rect 361842 130294 361898 130350
rect 361718 130170 361774 130226
rect 361842 130170 361898 130226
rect 361718 130046 361774 130102
rect 361842 130046 361898 130102
rect 361718 129922 361774 129978
rect 361842 129922 361898 129978
rect 392438 130294 392494 130350
rect 392562 130294 392618 130350
rect 392438 130170 392494 130226
rect 392562 130170 392618 130226
rect 392438 130046 392494 130102
rect 392562 130046 392618 130102
rect 392438 129922 392494 129978
rect 392562 129922 392618 129978
rect 423158 130294 423214 130350
rect 423282 130294 423338 130350
rect 423158 130170 423214 130226
rect 423282 130170 423338 130226
rect 423158 130046 423214 130102
rect 423282 130046 423338 130102
rect 423158 129922 423214 129978
rect 423282 129922 423338 129978
rect 453878 130294 453934 130350
rect 454002 130294 454058 130350
rect 453878 130170 453934 130226
rect 454002 130170 454058 130226
rect 453878 130046 453934 130102
rect 454002 130046 454058 130102
rect 453878 129922 453934 129978
rect 454002 129922 454058 129978
rect 484598 130294 484654 130350
rect 484722 130294 484778 130350
rect 484598 130170 484654 130226
rect 484722 130170 484778 130226
rect 484598 130046 484654 130102
rect 484722 130046 484778 130102
rect 484598 129922 484654 129978
rect 484722 129922 484778 129978
rect 515318 130294 515374 130350
rect 515442 130294 515498 130350
rect 515318 130170 515374 130226
rect 515442 130170 515498 130226
rect 515318 130046 515374 130102
rect 515442 130046 515498 130102
rect 515318 129922 515374 129978
rect 515442 129922 515498 129978
rect 546038 130294 546094 130350
rect 546162 130294 546218 130350
rect 546038 130170 546094 130226
rect 546162 130170 546218 130226
rect 546038 130046 546094 130102
rect 546162 130046 546218 130102
rect 546038 129922 546094 129978
rect 546162 129922 546218 129978
rect 561250 130294 561306 130350
rect 561374 130294 561430 130350
rect 561498 130294 561554 130350
rect 561622 130294 561678 130350
rect 561250 130170 561306 130226
rect 561374 130170 561430 130226
rect 561498 130170 561554 130226
rect 561622 130170 561678 130226
rect 561250 130046 561306 130102
rect 561374 130046 561430 130102
rect 561498 130046 561554 130102
rect 561622 130046 561678 130102
rect 561250 129922 561306 129978
rect 561374 129922 561430 129978
rect 561498 129922 561554 129978
rect 561622 129922 561678 129978
rect 131318 118294 131374 118350
rect 131442 118294 131498 118350
rect 131318 118170 131374 118226
rect 131442 118170 131498 118226
rect 131318 118046 131374 118102
rect 131442 118046 131498 118102
rect 131318 117922 131374 117978
rect 131442 117922 131498 117978
rect 162038 118294 162094 118350
rect 162162 118294 162218 118350
rect 162038 118170 162094 118226
rect 162162 118170 162218 118226
rect 162038 118046 162094 118102
rect 162162 118046 162218 118102
rect 162038 117922 162094 117978
rect 162162 117922 162218 117978
rect 192758 118294 192814 118350
rect 192882 118294 192938 118350
rect 192758 118170 192814 118226
rect 192882 118170 192938 118226
rect 192758 118046 192814 118102
rect 192882 118046 192938 118102
rect 192758 117922 192814 117978
rect 192882 117922 192938 117978
rect 223478 118294 223534 118350
rect 223602 118294 223658 118350
rect 223478 118170 223534 118226
rect 223602 118170 223658 118226
rect 223478 118046 223534 118102
rect 223602 118046 223658 118102
rect 223478 117922 223534 117978
rect 223602 117922 223658 117978
rect 254198 118294 254254 118350
rect 254322 118294 254378 118350
rect 254198 118170 254254 118226
rect 254322 118170 254378 118226
rect 254198 118046 254254 118102
rect 254322 118046 254378 118102
rect 254198 117922 254254 117978
rect 254322 117922 254378 117978
rect 284918 118294 284974 118350
rect 285042 118294 285098 118350
rect 284918 118170 284974 118226
rect 285042 118170 285098 118226
rect 284918 118046 284974 118102
rect 285042 118046 285098 118102
rect 284918 117922 284974 117978
rect 285042 117922 285098 117978
rect 315638 118294 315694 118350
rect 315762 118294 315818 118350
rect 315638 118170 315694 118226
rect 315762 118170 315818 118226
rect 315638 118046 315694 118102
rect 315762 118046 315818 118102
rect 315638 117922 315694 117978
rect 315762 117922 315818 117978
rect 346358 118294 346414 118350
rect 346482 118294 346538 118350
rect 346358 118170 346414 118226
rect 346482 118170 346538 118226
rect 346358 118046 346414 118102
rect 346482 118046 346538 118102
rect 346358 117922 346414 117978
rect 346482 117922 346538 117978
rect 377078 118294 377134 118350
rect 377202 118294 377258 118350
rect 377078 118170 377134 118226
rect 377202 118170 377258 118226
rect 377078 118046 377134 118102
rect 377202 118046 377258 118102
rect 377078 117922 377134 117978
rect 377202 117922 377258 117978
rect 407798 118294 407854 118350
rect 407922 118294 407978 118350
rect 407798 118170 407854 118226
rect 407922 118170 407978 118226
rect 407798 118046 407854 118102
rect 407922 118046 407978 118102
rect 407798 117922 407854 117978
rect 407922 117922 407978 117978
rect 438518 118294 438574 118350
rect 438642 118294 438698 118350
rect 438518 118170 438574 118226
rect 438642 118170 438698 118226
rect 438518 118046 438574 118102
rect 438642 118046 438698 118102
rect 438518 117922 438574 117978
rect 438642 117922 438698 117978
rect 469238 118294 469294 118350
rect 469362 118294 469418 118350
rect 469238 118170 469294 118226
rect 469362 118170 469418 118226
rect 469238 118046 469294 118102
rect 469362 118046 469418 118102
rect 469238 117922 469294 117978
rect 469362 117922 469418 117978
rect 499958 118294 500014 118350
rect 500082 118294 500138 118350
rect 499958 118170 500014 118226
rect 500082 118170 500138 118226
rect 499958 118046 500014 118102
rect 500082 118046 500138 118102
rect 499958 117922 500014 117978
rect 500082 117922 500138 117978
rect 530678 118294 530734 118350
rect 530802 118294 530858 118350
rect 530678 118170 530734 118226
rect 530802 118170 530858 118226
rect 530678 118046 530734 118102
rect 530802 118046 530858 118102
rect 530678 117922 530734 117978
rect 530802 117922 530858 117978
rect 111250 112294 111306 112350
rect 111374 112294 111430 112350
rect 111498 112294 111554 112350
rect 111622 112294 111678 112350
rect 111250 112170 111306 112226
rect 111374 112170 111430 112226
rect 111498 112170 111554 112226
rect 111622 112170 111678 112226
rect 111250 112046 111306 112102
rect 111374 112046 111430 112102
rect 111498 112046 111554 112102
rect 111622 112046 111678 112102
rect 111250 111922 111306 111978
rect 111374 111922 111430 111978
rect 111498 111922 111554 111978
rect 111622 111922 111678 111978
rect 96970 100294 97026 100350
rect 97094 100294 97150 100350
rect 97218 100294 97274 100350
rect 97342 100294 97398 100350
rect 96970 100170 97026 100226
rect 97094 100170 97150 100226
rect 97218 100170 97274 100226
rect 97342 100170 97398 100226
rect 96970 100046 97026 100102
rect 97094 100046 97150 100102
rect 97218 100046 97274 100102
rect 97342 100046 97398 100102
rect 96970 99922 97026 99978
rect 97094 99922 97150 99978
rect 97218 99922 97274 99978
rect 97342 99922 97398 99978
rect 100598 100294 100654 100350
rect 100722 100294 100778 100350
rect 100598 100170 100654 100226
rect 100722 100170 100778 100226
rect 100598 100046 100654 100102
rect 100722 100046 100778 100102
rect 100598 99922 100654 99978
rect 100722 99922 100778 99978
rect 115958 112294 116014 112350
rect 116082 112294 116138 112350
rect 115958 112170 116014 112226
rect 116082 112170 116138 112226
rect 115958 112046 116014 112102
rect 116082 112046 116138 112102
rect 115958 111922 116014 111978
rect 116082 111922 116138 111978
rect 146678 112294 146734 112350
rect 146802 112294 146858 112350
rect 146678 112170 146734 112226
rect 146802 112170 146858 112226
rect 146678 112046 146734 112102
rect 146802 112046 146858 112102
rect 146678 111922 146734 111978
rect 146802 111922 146858 111978
rect 177398 112294 177454 112350
rect 177522 112294 177578 112350
rect 177398 112170 177454 112226
rect 177522 112170 177578 112226
rect 177398 112046 177454 112102
rect 177522 112046 177578 112102
rect 177398 111922 177454 111978
rect 177522 111922 177578 111978
rect 208118 112294 208174 112350
rect 208242 112294 208298 112350
rect 208118 112170 208174 112226
rect 208242 112170 208298 112226
rect 208118 112046 208174 112102
rect 208242 112046 208298 112102
rect 208118 111922 208174 111978
rect 208242 111922 208298 111978
rect 238838 112294 238894 112350
rect 238962 112294 239018 112350
rect 238838 112170 238894 112226
rect 238962 112170 239018 112226
rect 238838 112046 238894 112102
rect 238962 112046 239018 112102
rect 238838 111922 238894 111978
rect 238962 111922 239018 111978
rect 269558 112294 269614 112350
rect 269682 112294 269738 112350
rect 269558 112170 269614 112226
rect 269682 112170 269738 112226
rect 269558 112046 269614 112102
rect 269682 112046 269738 112102
rect 269558 111922 269614 111978
rect 269682 111922 269738 111978
rect 300278 112294 300334 112350
rect 300402 112294 300458 112350
rect 300278 112170 300334 112226
rect 300402 112170 300458 112226
rect 300278 112046 300334 112102
rect 300402 112046 300458 112102
rect 300278 111922 300334 111978
rect 300402 111922 300458 111978
rect 330998 112294 331054 112350
rect 331122 112294 331178 112350
rect 330998 112170 331054 112226
rect 331122 112170 331178 112226
rect 330998 112046 331054 112102
rect 331122 112046 331178 112102
rect 330998 111922 331054 111978
rect 331122 111922 331178 111978
rect 361718 112294 361774 112350
rect 361842 112294 361898 112350
rect 361718 112170 361774 112226
rect 361842 112170 361898 112226
rect 361718 112046 361774 112102
rect 361842 112046 361898 112102
rect 361718 111922 361774 111978
rect 361842 111922 361898 111978
rect 392438 112294 392494 112350
rect 392562 112294 392618 112350
rect 392438 112170 392494 112226
rect 392562 112170 392618 112226
rect 392438 112046 392494 112102
rect 392562 112046 392618 112102
rect 392438 111922 392494 111978
rect 392562 111922 392618 111978
rect 423158 112294 423214 112350
rect 423282 112294 423338 112350
rect 423158 112170 423214 112226
rect 423282 112170 423338 112226
rect 423158 112046 423214 112102
rect 423282 112046 423338 112102
rect 423158 111922 423214 111978
rect 423282 111922 423338 111978
rect 453878 112294 453934 112350
rect 454002 112294 454058 112350
rect 453878 112170 453934 112226
rect 454002 112170 454058 112226
rect 453878 112046 453934 112102
rect 454002 112046 454058 112102
rect 453878 111922 453934 111978
rect 454002 111922 454058 111978
rect 484598 112294 484654 112350
rect 484722 112294 484778 112350
rect 484598 112170 484654 112226
rect 484722 112170 484778 112226
rect 484598 112046 484654 112102
rect 484722 112046 484778 112102
rect 484598 111922 484654 111978
rect 484722 111922 484778 111978
rect 515318 112294 515374 112350
rect 515442 112294 515498 112350
rect 515318 112170 515374 112226
rect 515442 112170 515498 112226
rect 515318 112046 515374 112102
rect 515442 112046 515498 112102
rect 515318 111922 515374 111978
rect 515442 111922 515498 111978
rect 546038 112294 546094 112350
rect 546162 112294 546218 112350
rect 546038 112170 546094 112226
rect 546162 112170 546218 112226
rect 546038 112046 546094 112102
rect 546162 112046 546218 112102
rect 546038 111922 546094 111978
rect 546162 111922 546218 111978
rect 561250 112294 561306 112350
rect 561374 112294 561430 112350
rect 561498 112294 561554 112350
rect 561622 112294 561678 112350
rect 561250 112170 561306 112226
rect 561374 112170 561430 112226
rect 561498 112170 561554 112226
rect 561622 112170 561678 112226
rect 561250 112046 561306 112102
rect 561374 112046 561430 112102
rect 561498 112046 561554 112102
rect 561622 112046 561678 112102
rect 561250 111922 561306 111978
rect 561374 111922 561430 111978
rect 561498 111922 561554 111978
rect 561622 111922 561678 111978
rect 131318 100294 131374 100350
rect 131442 100294 131498 100350
rect 131318 100170 131374 100226
rect 131442 100170 131498 100226
rect 131318 100046 131374 100102
rect 131442 100046 131498 100102
rect 131318 99922 131374 99978
rect 131442 99922 131498 99978
rect 162038 100294 162094 100350
rect 162162 100294 162218 100350
rect 162038 100170 162094 100226
rect 162162 100170 162218 100226
rect 162038 100046 162094 100102
rect 162162 100046 162218 100102
rect 162038 99922 162094 99978
rect 162162 99922 162218 99978
rect 192758 100294 192814 100350
rect 192882 100294 192938 100350
rect 192758 100170 192814 100226
rect 192882 100170 192938 100226
rect 192758 100046 192814 100102
rect 192882 100046 192938 100102
rect 192758 99922 192814 99978
rect 192882 99922 192938 99978
rect 223478 100294 223534 100350
rect 223602 100294 223658 100350
rect 223478 100170 223534 100226
rect 223602 100170 223658 100226
rect 223478 100046 223534 100102
rect 223602 100046 223658 100102
rect 223478 99922 223534 99978
rect 223602 99922 223658 99978
rect 254198 100294 254254 100350
rect 254322 100294 254378 100350
rect 254198 100170 254254 100226
rect 254322 100170 254378 100226
rect 254198 100046 254254 100102
rect 254322 100046 254378 100102
rect 254198 99922 254254 99978
rect 254322 99922 254378 99978
rect 284918 100294 284974 100350
rect 285042 100294 285098 100350
rect 284918 100170 284974 100226
rect 285042 100170 285098 100226
rect 284918 100046 284974 100102
rect 285042 100046 285098 100102
rect 284918 99922 284974 99978
rect 285042 99922 285098 99978
rect 315638 100294 315694 100350
rect 315762 100294 315818 100350
rect 315638 100170 315694 100226
rect 315762 100170 315818 100226
rect 315638 100046 315694 100102
rect 315762 100046 315818 100102
rect 315638 99922 315694 99978
rect 315762 99922 315818 99978
rect 346358 100294 346414 100350
rect 346482 100294 346538 100350
rect 346358 100170 346414 100226
rect 346482 100170 346538 100226
rect 346358 100046 346414 100102
rect 346482 100046 346538 100102
rect 346358 99922 346414 99978
rect 346482 99922 346538 99978
rect 377078 100294 377134 100350
rect 377202 100294 377258 100350
rect 377078 100170 377134 100226
rect 377202 100170 377258 100226
rect 377078 100046 377134 100102
rect 377202 100046 377258 100102
rect 377078 99922 377134 99978
rect 377202 99922 377258 99978
rect 407798 100294 407854 100350
rect 407922 100294 407978 100350
rect 407798 100170 407854 100226
rect 407922 100170 407978 100226
rect 407798 100046 407854 100102
rect 407922 100046 407978 100102
rect 407798 99922 407854 99978
rect 407922 99922 407978 99978
rect 438518 100294 438574 100350
rect 438642 100294 438698 100350
rect 438518 100170 438574 100226
rect 438642 100170 438698 100226
rect 438518 100046 438574 100102
rect 438642 100046 438698 100102
rect 438518 99922 438574 99978
rect 438642 99922 438698 99978
rect 469238 100294 469294 100350
rect 469362 100294 469418 100350
rect 469238 100170 469294 100226
rect 469362 100170 469418 100226
rect 469238 100046 469294 100102
rect 469362 100046 469418 100102
rect 469238 99922 469294 99978
rect 469362 99922 469418 99978
rect 499958 100294 500014 100350
rect 500082 100294 500138 100350
rect 499958 100170 500014 100226
rect 500082 100170 500138 100226
rect 499958 100046 500014 100102
rect 500082 100046 500138 100102
rect 499958 99922 500014 99978
rect 500082 99922 500138 99978
rect 530678 100294 530734 100350
rect 530802 100294 530858 100350
rect 530678 100170 530734 100226
rect 530802 100170 530858 100226
rect 530678 100046 530734 100102
rect 530802 100046 530858 100102
rect 530678 99922 530734 99978
rect 530802 99922 530858 99978
rect 111250 94294 111306 94350
rect 111374 94294 111430 94350
rect 111498 94294 111554 94350
rect 111622 94294 111678 94350
rect 111250 94170 111306 94226
rect 111374 94170 111430 94226
rect 111498 94170 111554 94226
rect 111622 94170 111678 94226
rect 111250 94046 111306 94102
rect 111374 94046 111430 94102
rect 111498 94046 111554 94102
rect 111622 94046 111678 94102
rect 111250 93922 111306 93978
rect 111374 93922 111430 93978
rect 111498 93922 111554 93978
rect 111622 93922 111678 93978
rect 96970 82294 97026 82350
rect 97094 82294 97150 82350
rect 97218 82294 97274 82350
rect 97342 82294 97398 82350
rect 96970 82170 97026 82226
rect 97094 82170 97150 82226
rect 97218 82170 97274 82226
rect 97342 82170 97398 82226
rect 96970 82046 97026 82102
rect 97094 82046 97150 82102
rect 97218 82046 97274 82102
rect 97342 82046 97398 82102
rect 96970 81922 97026 81978
rect 97094 81922 97150 81978
rect 97218 81922 97274 81978
rect 97342 81922 97398 81978
rect 100598 82294 100654 82350
rect 100722 82294 100778 82350
rect 100598 82170 100654 82226
rect 100722 82170 100778 82226
rect 100598 82046 100654 82102
rect 100722 82046 100778 82102
rect 100598 81922 100654 81978
rect 100722 81922 100778 81978
rect 115958 94294 116014 94350
rect 116082 94294 116138 94350
rect 115958 94170 116014 94226
rect 116082 94170 116138 94226
rect 115958 94046 116014 94102
rect 116082 94046 116138 94102
rect 115958 93922 116014 93978
rect 116082 93922 116138 93978
rect 146678 94294 146734 94350
rect 146802 94294 146858 94350
rect 146678 94170 146734 94226
rect 146802 94170 146858 94226
rect 146678 94046 146734 94102
rect 146802 94046 146858 94102
rect 146678 93922 146734 93978
rect 146802 93922 146858 93978
rect 177398 94294 177454 94350
rect 177522 94294 177578 94350
rect 177398 94170 177454 94226
rect 177522 94170 177578 94226
rect 177398 94046 177454 94102
rect 177522 94046 177578 94102
rect 177398 93922 177454 93978
rect 177522 93922 177578 93978
rect 208118 94294 208174 94350
rect 208242 94294 208298 94350
rect 208118 94170 208174 94226
rect 208242 94170 208298 94226
rect 208118 94046 208174 94102
rect 208242 94046 208298 94102
rect 208118 93922 208174 93978
rect 208242 93922 208298 93978
rect 238838 94294 238894 94350
rect 238962 94294 239018 94350
rect 238838 94170 238894 94226
rect 238962 94170 239018 94226
rect 238838 94046 238894 94102
rect 238962 94046 239018 94102
rect 238838 93922 238894 93978
rect 238962 93922 239018 93978
rect 269558 94294 269614 94350
rect 269682 94294 269738 94350
rect 269558 94170 269614 94226
rect 269682 94170 269738 94226
rect 269558 94046 269614 94102
rect 269682 94046 269738 94102
rect 269558 93922 269614 93978
rect 269682 93922 269738 93978
rect 300278 94294 300334 94350
rect 300402 94294 300458 94350
rect 300278 94170 300334 94226
rect 300402 94170 300458 94226
rect 300278 94046 300334 94102
rect 300402 94046 300458 94102
rect 300278 93922 300334 93978
rect 300402 93922 300458 93978
rect 330998 94294 331054 94350
rect 331122 94294 331178 94350
rect 330998 94170 331054 94226
rect 331122 94170 331178 94226
rect 330998 94046 331054 94102
rect 331122 94046 331178 94102
rect 330998 93922 331054 93978
rect 331122 93922 331178 93978
rect 361718 94294 361774 94350
rect 361842 94294 361898 94350
rect 361718 94170 361774 94226
rect 361842 94170 361898 94226
rect 361718 94046 361774 94102
rect 361842 94046 361898 94102
rect 361718 93922 361774 93978
rect 361842 93922 361898 93978
rect 392438 94294 392494 94350
rect 392562 94294 392618 94350
rect 392438 94170 392494 94226
rect 392562 94170 392618 94226
rect 392438 94046 392494 94102
rect 392562 94046 392618 94102
rect 392438 93922 392494 93978
rect 392562 93922 392618 93978
rect 423158 94294 423214 94350
rect 423282 94294 423338 94350
rect 423158 94170 423214 94226
rect 423282 94170 423338 94226
rect 423158 94046 423214 94102
rect 423282 94046 423338 94102
rect 423158 93922 423214 93978
rect 423282 93922 423338 93978
rect 453878 94294 453934 94350
rect 454002 94294 454058 94350
rect 453878 94170 453934 94226
rect 454002 94170 454058 94226
rect 453878 94046 453934 94102
rect 454002 94046 454058 94102
rect 453878 93922 453934 93978
rect 454002 93922 454058 93978
rect 484598 94294 484654 94350
rect 484722 94294 484778 94350
rect 484598 94170 484654 94226
rect 484722 94170 484778 94226
rect 484598 94046 484654 94102
rect 484722 94046 484778 94102
rect 484598 93922 484654 93978
rect 484722 93922 484778 93978
rect 515318 94294 515374 94350
rect 515442 94294 515498 94350
rect 515318 94170 515374 94226
rect 515442 94170 515498 94226
rect 515318 94046 515374 94102
rect 515442 94046 515498 94102
rect 515318 93922 515374 93978
rect 515442 93922 515498 93978
rect 546038 94294 546094 94350
rect 546162 94294 546218 94350
rect 546038 94170 546094 94226
rect 546162 94170 546218 94226
rect 546038 94046 546094 94102
rect 546162 94046 546218 94102
rect 546038 93922 546094 93978
rect 546162 93922 546218 93978
rect 561250 94294 561306 94350
rect 561374 94294 561430 94350
rect 561498 94294 561554 94350
rect 561622 94294 561678 94350
rect 561250 94170 561306 94226
rect 561374 94170 561430 94226
rect 561498 94170 561554 94226
rect 561622 94170 561678 94226
rect 561250 94046 561306 94102
rect 561374 94046 561430 94102
rect 561498 94046 561554 94102
rect 561622 94046 561678 94102
rect 561250 93922 561306 93978
rect 561374 93922 561430 93978
rect 561498 93922 561554 93978
rect 561622 93922 561678 93978
rect 131318 82294 131374 82350
rect 131442 82294 131498 82350
rect 131318 82170 131374 82226
rect 131442 82170 131498 82226
rect 131318 82046 131374 82102
rect 131442 82046 131498 82102
rect 131318 81922 131374 81978
rect 131442 81922 131498 81978
rect 162038 82294 162094 82350
rect 162162 82294 162218 82350
rect 162038 82170 162094 82226
rect 162162 82170 162218 82226
rect 162038 82046 162094 82102
rect 162162 82046 162218 82102
rect 162038 81922 162094 81978
rect 162162 81922 162218 81978
rect 192758 82294 192814 82350
rect 192882 82294 192938 82350
rect 192758 82170 192814 82226
rect 192882 82170 192938 82226
rect 192758 82046 192814 82102
rect 192882 82046 192938 82102
rect 192758 81922 192814 81978
rect 192882 81922 192938 81978
rect 223478 82294 223534 82350
rect 223602 82294 223658 82350
rect 223478 82170 223534 82226
rect 223602 82170 223658 82226
rect 223478 82046 223534 82102
rect 223602 82046 223658 82102
rect 223478 81922 223534 81978
rect 223602 81922 223658 81978
rect 254198 82294 254254 82350
rect 254322 82294 254378 82350
rect 254198 82170 254254 82226
rect 254322 82170 254378 82226
rect 254198 82046 254254 82102
rect 254322 82046 254378 82102
rect 254198 81922 254254 81978
rect 254322 81922 254378 81978
rect 284918 82294 284974 82350
rect 285042 82294 285098 82350
rect 284918 82170 284974 82226
rect 285042 82170 285098 82226
rect 284918 82046 284974 82102
rect 285042 82046 285098 82102
rect 284918 81922 284974 81978
rect 285042 81922 285098 81978
rect 315638 82294 315694 82350
rect 315762 82294 315818 82350
rect 315638 82170 315694 82226
rect 315762 82170 315818 82226
rect 315638 82046 315694 82102
rect 315762 82046 315818 82102
rect 315638 81922 315694 81978
rect 315762 81922 315818 81978
rect 346358 82294 346414 82350
rect 346482 82294 346538 82350
rect 346358 82170 346414 82226
rect 346482 82170 346538 82226
rect 346358 82046 346414 82102
rect 346482 82046 346538 82102
rect 346358 81922 346414 81978
rect 346482 81922 346538 81978
rect 377078 82294 377134 82350
rect 377202 82294 377258 82350
rect 377078 82170 377134 82226
rect 377202 82170 377258 82226
rect 377078 82046 377134 82102
rect 377202 82046 377258 82102
rect 377078 81922 377134 81978
rect 377202 81922 377258 81978
rect 407798 82294 407854 82350
rect 407922 82294 407978 82350
rect 407798 82170 407854 82226
rect 407922 82170 407978 82226
rect 407798 82046 407854 82102
rect 407922 82046 407978 82102
rect 407798 81922 407854 81978
rect 407922 81922 407978 81978
rect 438518 82294 438574 82350
rect 438642 82294 438698 82350
rect 438518 82170 438574 82226
rect 438642 82170 438698 82226
rect 438518 82046 438574 82102
rect 438642 82046 438698 82102
rect 438518 81922 438574 81978
rect 438642 81922 438698 81978
rect 469238 82294 469294 82350
rect 469362 82294 469418 82350
rect 469238 82170 469294 82226
rect 469362 82170 469418 82226
rect 469238 82046 469294 82102
rect 469362 82046 469418 82102
rect 469238 81922 469294 81978
rect 469362 81922 469418 81978
rect 499958 82294 500014 82350
rect 500082 82294 500138 82350
rect 499958 82170 500014 82226
rect 500082 82170 500138 82226
rect 499958 82046 500014 82102
rect 500082 82046 500138 82102
rect 499958 81922 500014 81978
rect 500082 81922 500138 81978
rect 530678 82294 530734 82350
rect 530802 82294 530858 82350
rect 530678 82170 530734 82226
rect 530802 82170 530858 82226
rect 530678 82046 530734 82102
rect 530802 82046 530858 82102
rect 530678 81922 530734 81978
rect 530802 81922 530858 81978
rect 111250 76294 111306 76350
rect 111374 76294 111430 76350
rect 111498 76294 111554 76350
rect 111622 76294 111678 76350
rect 111250 76170 111306 76226
rect 111374 76170 111430 76226
rect 111498 76170 111554 76226
rect 111622 76170 111678 76226
rect 111250 76046 111306 76102
rect 111374 76046 111430 76102
rect 111498 76046 111554 76102
rect 111622 76046 111678 76102
rect 111250 75922 111306 75978
rect 111374 75922 111430 75978
rect 111498 75922 111554 75978
rect 111622 75922 111678 75978
rect 96970 64294 97026 64350
rect 97094 64294 97150 64350
rect 97218 64294 97274 64350
rect 97342 64294 97398 64350
rect 96970 64170 97026 64226
rect 97094 64170 97150 64226
rect 97218 64170 97274 64226
rect 97342 64170 97398 64226
rect 96970 64046 97026 64102
rect 97094 64046 97150 64102
rect 97218 64046 97274 64102
rect 97342 64046 97398 64102
rect 96970 63922 97026 63978
rect 97094 63922 97150 63978
rect 97218 63922 97274 63978
rect 97342 63922 97398 63978
rect 100598 64294 100654 64350
rect 100722 64294 100778 64350
rect 100598 64170 100654 64226
rect 100722 64170 100778 64226
rect 100598 64046 100654 64102
rect 100722 64046 100778 64102
rect 100598 63922 100654 63978
rect 100722 63922 100778 63978
rect 115958 76294 116014 76350
rect 116082 76294 116138 76350
rect 115958 76170 116014 76226
rect 116082 76170 116138 76226
rect 115958 76046 116014 76102
rect 116082 76046 116138 76102
rect 115958 75922 116014 75978
rect 116082 75922 116138 75978
rect 146678 76294 146734 76350
rect 146802 76294 146858 76350
rect 146678 76170 146734 76226
rect 146802 76170 146858 76226
rect 146678 76046 146734 76102
rect 146802 76046 146858 76102
rect 146678 75922 146734 75978
rect 146802 75922 146858 75978
rect 177398 76294 177454 76350
rect 177522 76294 177578 76350
rect 177398 76170 177454 76226
rect 177522 76170 177578 76226
rect 177398 76046 177454 76102
rect 177522 76046 177578 76102
rect 177398 75922 177454 75978
rect 177522 75922 177578 75978
rect 208118 76294 208174 76350
rect 208242 76294 208298 76350
rect 208118 76170 208174 76226
rect 208242 76170 208298 76226
rect 208118 76046 208174 76102
rect 208242 76046 208298 76102
rect 208118 75922 208174 75978
rect 208242 75922 208298 75978
rect 238838 76294 238894 76350
rect 238962 76294 239018 76350
rect 238838 76170 238894 76226
rect 238962 76170 239018 76226
rect 238838 76046 238894 76102
rect 238962 76046 239018 76102
rect 238838 75922 238894 75978
rect 238962 75922 239018 75978
rect 269558 76294 269614 76350
rect 269682 76294 269738 76350
rect 269558 76170 269614 76226
rect 269682 76170 269738 76226
rect 269558 76046 269614 76102
rect 269682 76046 269738 76102
rect 269558 75922 269614 75978
rect 269682 75922 269738 75978
rect 300278 76294 300334 76350
rect 300402 76294 300458 76350
rect 300278 76170 300334 76226
rect 300402 76170 300458 76226
rect 300278 76046 300334 76102
rect 300402 76046 300458 76102
rect 300278 75922 300334 75978
rect 300402 75922 300458 75978
rect 330998 76294 331054 76350
rect 331122 76294 331178 76350
rect 330998 76170 331054 76226
rect 331122 76170 331178 76226
rect 330998 76046 331054 76102
rect 331122 76046 331178 76102
rect 330998 75922 331054 75978
rect 331122 75922 331178 75978
rect 361718 76294 361774 76350
rect 361842 76294 361898 76350
rect 361718 76170 361774 76226
rect 361842 76170 361898 76226
rect 361718 76046 361774 76102
rect 361842 76046 361898 76102
rect 361718 75922 361774 75978
rect 361842 75922 361898 75978
rect 392438 76294 392494 76350
rect 392562 76294 392618 76350
rect 392438 76170 392494 76226
rect 392562 76170 392618 76226
rect 392438 76046 392494 76102
rect 392562 76046 392618 76102
rect 392438 75922 392494 75978
rect 392562 75922 392618 75978
rect 423158 76294 423214 76350
rect 423282 76294 423338 76350
rect 423158 76170 423214 76226
rect 423282 76170 423338 76226
rect 423158 76046 423214 76102
rect 423282 76046 423338 76102
rect 423158 75922 423214 75978
rect 423282 75922 423338 75978
rect 453878 76294 453934 76350
rect 454002 76294 454058 76350
rect 453878 76170 453934 76226
rect 454002 76170 454058 76226
rect 453878 76046 453934 76102
rect 454002 76046 454058 76102
rect 453878 75922 453934 75978
rect 454002 75922 454058 75978
rect 484598 76294 484654 76350
rect 484722 76294 484778 76350
rect 484598 76170 484654 76226
rect 484722 76170 484778 76226
rect 484598 76046 484654 76102
rect 484722 76046 484778 76102
rect 484598 75922 484654 75978
rect 484722 75922 484778 75978
rect 515318 76294 515374 76350
rect 515442 76294 515498 76350
rect 515318 76170 515374 76226
rect 515442 76170 515498 76226
rect 515318 76046 515374 76102
rect 515442 76046 515498 76102
rect 515318 75922 515374 75978
rect 515442 75922 515498 75978
rect 546038 76294 546094 76350
rect 546162 76294 546218 76350
rect 546038 76170 546094 76226
rect 546162 76170 546218 76226
rect 546038 76046 546094 76102
rect 546162 76046 546218 76102
rect 546038 75922 546094 75978
rect 546162 75922 546218 75978
rect 561250 76294 561306 76350
rect 561374 76294 561430 76350
rect 561498 76294 561554 76350
rect 561622 76294 561678 76350
rect 561250 76170 561306 76226
rect 561374 76170 561430 76226
rect 561498 76170 561554 76226
rect 561622 76170 561678 76226
rect 561250 76046 561306 76102
rect 561374 76046 561430 76102
rect 561498 76046 561554 76102
rect 561622 76046 561678 76102
rect 561250 75922 561306 75978
rect 561374 75922 561430 75978
rect 561498 75922 561554 75978
rect 561622 75922 561678 75978
rect 131318 64294 131374 64350
rect 131442 64294 131498 64350
rect 131318 64170 131374 64226
rect 131442 64170 131498 64226
rect 131318 64046 131374 64102
rect 131442 64046 131498 64102
rect 131318 63922 131374 63978
rect 131442 63922 131498 63978
rect 162038 64294 162094 64350
rect 162162 64294 162218 64350
rect 162038 64170 162094 64226
rect 162162 64170 162218 64226
rect 162038 64046 162094 64102
rect 162162 64046 162218 64102
rect 162038 63922 162094 63978
rect 162162 63922 162218 63978
rect 192758 64294 192814 64350
rect 192882 64294 192938 64350
rect 192758 64170 192814 64226
rect 192882 64170 192938 64226
rect 192758 64046 192814 64102
rect 192882 64046 192938 64102
rect 192758 63922 192814 63978
rect 192882 63922 192938 63978
rect 223478 64294 223534 64350
rect 223602 64294 223658 64350
rect 223478 64170 223534 64226
rect 223602 64170 223658 64226
rect 223478 64046 223534 64102
rect 223602 64046 223658 64102
rect 223478 63922 223534 63978
rect 223602 63922 223658 63978
rect 254198 64294 254254 64350
rect 254322 64294 254378 64350
rect 254198 64170 254254 64226
rect 254322 64170 254378 64226
rect 254198 64046 254254 64102
rect 254322 64046 254378 64102
rect 254198 63922 254254 63978
rect 254322 63922 254378 63978
rect 284918 64294 284974 64350
rect 285042 64294 285098 64350
rect 284918 64170 284974 64226
rect 285042 64170 285098 64226
rect 284918 64046 284974 64102
rect 285042 64046 285098 64102
rect 284918 63922 284974 63978
rect 285042 63922 285098 63978
rect 315638 64294 315694 64350
rect 315762 64294 315818 64350
rect 315638 64170 315694 64226
rect 315762 64170 315818 64226
rect 315638 64046 315694 64102
rect 315762 64046 315818 64102
rect 315638 63922 315694 63978
rect 315762 63922 315818 63978
rect 346358 64294 346414 64350
rect 346482 64294 346538 64350
rect 346358 64170 346414 64226
rect 346482 64170 346538 64226
rect 346358 64046 346414 64102
rect 346482 64046 346538 64102
rect 346358 63922 346414 63978
rect 346482 63922 346538 63978
rect 377078 64294 377134 64350
rect 377202 64294 377258 64350
rect 377078 64170 377134 64226
rect 377202 64170 377258 64226
rect 377078 64046 377134 64102
rect 377202 64046 377258 64102
rect 377078 63922 377134 63978
rect 377202 63922 377258 63978
rect 407798 64294 407854 64350
rect 407922 64294 407978 64350
rect 407798 64170 407854 64226
rect 407922 64170 407978 64226
rect 407798 64046 407854 64102
rect 407922 64046 407978 64102
rect 407798 63922 407854 63978
rect 407922 63922 407978 63978
rect 438518 64294 438574 64350
rect 438642 64294 438698 64350
rect 438518 64170 438574 64226
rect 438642 64170 438698 64226
rect 438518 64046 438574 64102
rect 438642 64046 438698 64102
rect 438518 63922 438574 63978
rect 438642 63922 438698 63978
rect 469238 64294 469294 64350
rect 469362 64294 469418 64350
rect 469238 64170 469294 64226
rect 469362 64170 469418 64226
rect 469238 64046 469294 64102
rect 469362 64046 469418 64102
rect 469238 63922 469294 63978
rect 469362 63922 469418 63978
rect 499958 64294 500014 64350
rect 500082 64294 500138 64350
rect 499958 64170 500014 64226
rect 500082 64170 500138 64226
rect 499958 64046 500014 64102
rect 500082 64046 500138 64102
rect 499958 63922 500014 63978
rect 500082 63922 500138 63978
rect 530678 64294 530734 64350
rect 530802 64294 530858 64350
rect 530678 64170 530734 64226
rect 530802 64170 530858 64226
rect 530678 64046 530734 64102
rect 530802 64046 530858 64102
rect 530678 63922 530734 63978
rect 530802 63922 530858 63978
rect 111250 58294 111306 58350
rect 111374 58294 111430 58350
rect 111498 58294 111554 58350
rect 111622 58294 111678 58350
rect 111250 58170 111306 58226
rect 111374 58170 111430 58226
rect 111498 58170 111554 58226
rect 111622 58170 111678 58226
rect 111250 58046 111306 58102
rect 111374 58046 111430 58102
rect 111498 58046 111554 58102
rect 111622 58046 111678 58102
rect 111250 57922 111306 57978
rect 111374 57922 111430 57978
rect 111498 57922 111554 57978
rect 111622 57922 111678 57978
rect 96970 46294 97026 46350
rect 97094 46294 97150 46350
rect 97218 46294 97274 46350
rect 97342 46294 97398 46350
rect 96970 46170 97026 46226
rect 97094 46170 97150 46226
rect 97218 46170 97274 46226
rect 97342 46170 97398 46226
rect 96970 46046 97026 46102
rect 97094 46046 97150 46102
rect 97218 46046 97274 46102
rect 97342 46046 97398 46102
rect 96970 45922 97026 45978
rect 97094 45922 97150 45978
rect 97218 45922 97274 45978
rect 97342 45922 97398 45978
rect 100598 46294 100654 46350
rect 100722 46294 100778 46350
rect 100598 46170 100654 46226
rect 100722 46170 100778 46226
rect 100598 46046 100654 46102
rect 100722 46046 100778 46102
rect 100598 45922 100654 45978
rect 100722 45922 100778 45978
rect 96970 28294 97026 28350
rect 97094 28294 97150 28350
rect 97218 28294 97274 28350
rect 97342 28294 97398 28350
rect 96970 28170 97026 28226
rect 97094 28170 97150 28226
rect 97218 28170 97274 28226
rect 97342 28170 97398 28226
rect 96970 28046 97026 28102
rect 97094 28046 97150 28102
rect 97218 28046 97274 28102
rect 97342 28046 97398 28102
rect 96970 27922 97026 27978
rect 97094 27922 97150 27978
rect 97218 27922 97274 27978
rect 97342 27922 97398 27978
rect 96970 10294 97026 10350
rect 97094 10294 97150 10350
rect 97218 10294 97274 10350
rect 97342 10294 97398 10350
rect 96970 10170 97026 10226
rect 97094 10170 97150 10226
rect 97218 10170 97274 10226
rect 97342 10170 97398 10226
rect 96970 10046 97026 10102
rect 97094 10046 97150 10102
rect 97218 10046 97274 10102
rect 97342 10046 97398 10102
rect 96970 9922 97026 9978
rect 97094 9922 97150 9978
rect 97218 9922 97274 9978
rect 97342 9922 97398 9978
rect 96970 -1176 97026 -1120
rect 97094 -1176 97150 -1120
rect 97218 -1176 97274 -1120
rect 97342 -1176 97398 -1120
rect 96970 -1300 97026 -1244
rect 97094 -1300 97150 -1244
rect 97218 -1300 97274 -1244
rect 97342 -1300 97398 -1244
rect 96970 -1424 97026 -1368
rect 97094 -1424 97150 -1368
rect 97218 -1424 97274 -1368
rect 97342 -1424 97398 -1368
rect 96970 -1548 97026 -1492
rect 97094 -1548 97150 -1492
rect 97218 -1548 97274 -1492
rect 97342 -1548 97398 -1492
rect 115958 58294 116014 58350
rect 116082 58294 116138 58350
rect 115958 58170 116014 58226
rect 116082 58170 116138 58226
rect 115958 58046 116014 58102
rect 116082 58046 116138 58102
rect 115958 57922 116014 57978
rect 116082 57922 116138 57978
rect 146678 58294 146734 58350
rect 146802 58294 146858 58350
rect 146678 58170 146734 58226
rect 146802 58170 146858 58226
rect 146678 58046 146734 58102
rect 146802 58046 146858 58102
rect 146678 57922 146734 57978
rect 146802 57922 146858 57978
rect 177398 58294 177454 58350
rect 177522 58294 177578 58350
rect 177398 58170 177454 58226
rect 177522 58170 177578 58226
rect 177398 58046 177454 58102
rect 177522 58046 177578 58102
rect 177398 57922 177454 57978
rect 177522 57922 177578 57978
rect 208118 58294 208174 58350
rect 208242 58294 208298 58350
rect 208118 58170 208174 58226
rect 208242 58170 208298 58226
rect 208118 58046 208174 58102
rect 208242 58046 208298 58102
rect 208118 57922 208174 57978
rect 208242 57922 208298 57978
rect 238838 58294 238894 58350
rect 238962 58294 239018 58350
rect 238838 58170 238894 58226
rect 238962 58170 239018 58226
rect 238838 58046 238894 58102
rect 238962 58046 239018 58102
rect 238838 57922 238894 57978
rect 238962 57922 239018 57978
rect 269558 58294 269614 58350
rect 269682 58294 269738 58350
rect 269558 58170 269614 58226
rect 269682 58170 269738 58226
rect 269558 58046 269614 58102
rect 269682 58046 269738 58102
rect 269558 57922 269614 57978
rect 269682 57922 269738 57978
rect 300278 58294 300334 58350
rect 300402 58294 300458 58350
rect 300278 58170 300334 58226
rect 300402 58170 300458 58226
rect 300278 58046 300334 58102
rect 300402 58046 300458 58102
rect 300278 57922 300334 57978
rect 300402 57922 300458 57978
rect 330998 58294 331054 58350
rect 331122 58294 331178 58350
rect 330998 58170 331054 58226
rect 331122 58170 331178 58226
rect 330998 58046 331054 58102
rect 331122 58046 331178 58102
rect 330998 57922 331054 57978
rect 331122 57922 331178 57978
rect 361718 58294 361774 58350
rect 361842 58294 361898 58350
rect 361718 58170 361774 58226
rect 361842 58170 361898 58226
rect 361718 58046 361774 58102
rect 361842 58046 361898 58102
rect 361718 57922 361774 57978
rect 361842 57922 361898 57978
rect 392438 58294 392494 58350
rect 392562 58294 392618 58350
rect 392438 58170 392494 58226
rect 392562 58170 392618 58226
rect 392438 58046 392494 58102
rect 392562 58046 392618 58102
rect 392438 57922 392494 57978
rect 392562 57922 392618 57978
rect 423158 58294 423214 58350
rect 423282 58294 423338 58350
rect 423158 58170 423214 58226
rect 423282 58170 423338 58226
rect 423158 58046 423214 58102
rect 423282 58046 423338 58102
rect 423158 57922 423214 57978
rect 423282 57922 423338 57978
rect 453878 58294 453934 58350
rect 454002 58294 454058 58350
rect 453878 58170 453934 58226
rect 454002 58170 454058 58226
rect 453878 58046 453934 58102
rect 454002 58046 454058 58102
rect 453878 57922 453934 57978
rect 454002 57922 454058 57978
rect 484598 58294 484654 58350
rect 484722 58294 484778 58350
rect 484598 58170 484654 58226
rect 484722 58170 484778 58226
rect 484598 58046 484654 58102
rect 484722 58046 484778 58102
rect 484598 57922 484654 57978
rect 484722 57922 484778 57978
rect 515318 58294 515374 58350
rect 515442 58294 515498 58350
rect 515318 58170 515374 58226
rect 515442 58170 515498 58226
rect 515318 58046 515374 58102
rect 515442 58046 515498 58102
rect 515318 57922 515374 57978
rect 515442 57922 515498 57978
rect 546038 58294 546094 58350
rect 546162 58294 546218 58350
rect 546038 58170 546094 58226
rect 546162 58170 546218 58226
rect 546038 58046 546094 58102
rect 546162 58046 546218 58102
rect 546038 57922 546094 57978
rect 546162 57922 546218 57978
rect 561250 58294 561306 58350
rect 561374 58294 561430 58350
rect 561498 58294 561554 58350
rect 561622 58294 561678 58350
rect 561250 58170 561306 58226
rect 561374 58170 561430 58226
rect 561498 58170 561554 58226
rect 561622 58170 561678 58226
rect 561250 58046 561306 58102
rect 561374 58046 561430 58102
rect 561498 58046 561554 58102
rect 561622 58046 561678 58102
rect 561250 57922 561306 57978
rect 561374 57922 561430 57978
rect 561498 57922 561554 57978
rect 561622 57922 561678 57978
rect 131318 46294 131374 46350
rect 131442 46294 131498 46350
rect 131318 46170 131374 46226
rect 131442 46170 131498 46226
rect 131318 46046 131374 46102
rect 131442 46046 131498 46102
rect 131318 45922 131374 45978
rect 131442 45922 131498 45978
rect 162038 46294 162094 46350
rect 162162 46294 162218 46350
rect 162038 46170 162094 46226
rect 162162 46170 162218 46226
rect 162038 46046 162094 46102
rect 162162 46046 162218 46102
rect 162038 45922 162094 45978
rect 162162 45922 162218 45978
rect 192758 46294 192814 46350
rect 192882 46294 192938 46350
rect 192758 46170 192814 46226
rect 192882 46170 192938 46226
rect 192758 46046 192814 46102
rect 192882 46046 192938 46102
rect 192758 45922 192814 45978
rect 192882 45922 192938 45978
rect 223478 46294 223534 46350
rect 223602 46294 223658 46350
rect 223478 46170 223534 46226
rect 223602 46170 223658 46226
rect 223478 46046 223534 46102
rect 223602 46046 223658 46102
rect 223478 45922 223534 45978
rect 223602 45922 223658 45978
rect 254198 46294 254254 46350
rect 254322 46294 254378 46350
rect 254198 46170 254254 46226
rect 254322 46170 254378 46226
rect 254198 46046 254254 46102
rect 254322 46046 254378 46102
rect 254198 45922 254254 45978
rect 254322 45922 254378 45978
rect 284918 46294 284974 46350
rect 285042 46294 285098 46350
rect 284918 46170 284974 46226
rect 285042 46170 285098 46226
rect 284918 46046 284974 46102
rect 285042 46046 285098 46102
rect 284918 45922 284974 45978
rect 285042 45922 285098 45978
rect 315638 46294 315694 46350
rect 315762 46294 315818 46350
rect 315638 46170 315694 46226
rect 315762 46170 315818 46226
rect 315638 46046 315694 46102
rect 315762 46046 315818 46102
rect 315638 45922 315694 45978
rect 315762 45922 315818 45978
rect 346358 46294 346414 46350
rect 346482 46294 346538 46350
rect 346358 46170 346414 46226
rect 346482 46170 346538 46226
rect 346358 46046 346414 46102
rect 346482 46046 346538 46102
rect 346358 45922 346414 45978
rect 346482 45922 346538 45978
rect 377078 46294 377134 46350
rect 377202 46294 377258 46350
rect 377078 46170 377134 46226
rect 377202 46170 377258 46226
rect 377078 46046 377134 46102
rect 377202 46046 377258 46102
rect 377078 45922 377134 45978
rect 377202 45922 377258 45978
rect 407798 46294 407854 46350
rect 407922 46294 407978 46350
rect 407798 46170 407854 46226
rect 407922 46170 407978 46226
rect 407798 46046 407854 46102
rect 407922 46046 407978 46102
rect 407798 45922 407854 45978
rect 407922 45922 407978 45978
rect 438518 46294 438574 46350
rect 438642 46294 438698 46350
rect 438518 46170 438574 46226
rect 438642 46170 438698 46226
rect 438518 46046 438574 46102
rect 438642 46046 438698 46102
rect 438518 45922 438574 45978
rect 438642 45922 438698 45978
rect 469238 46294 469294 46350
rect 469362 46294 469418 46350
rect 469238 46170 469294 46226
rect 469362 46170 469418 46226
rect 469238 46046 469294 46102
rect 469362 46046 469418 46102
rect 469238 45922 469294 45978
rect 469362 45922 469418 45978
rect 499958 46294 500014 46350
rect 500082 46294 500138 46350
rect 499958 46170 500014 46226
rect 500082 46170 500138 46226
rect 499958 46046 500014 46102
rect 500082 46046 500138 46102
rect 499958 45922 500014 45978
rect 500082 45922 500138 45978
rect 530678 46294 530734 46350
rect 530802 46294 530858 46350
rect 530678 46170 530734 46226
rect 530802 46170 530858 46226
rect 530678 46046 530734 46102
rect 530802 46046 530858 46102
rect 530678 45922 530734 45978
rect 530802 45922 530858 45978
rect 111250 40294 111306 40350
rect 111374 40294 111430 40350
rect 111498 40294 111554 40350
rect 111622 40294 111678 40350
rect 111250 40170 111306 40226
rect 111374 40170 111430 40226
rect 111498 40170 111554 40226
rect 111622 40170 111678 40226
rect 111250 40046 111306 40102
rect 111374 40046 111430 40102
rect 111498 40046 111554 40102
rect 111622 40046 111678 40102
rect 111250 39922 111306 39978
rect 111374 39922 111430 39978
rect 111498 39922 111554 39978
rect 111622 39922 111678 39978
rect 115958 40294 116014 40350
rect 116082 40294 116138 40350
rect 115958 40170 116014 40226
rect 116082 40170 116138 40226
rect 115958 40046 116014 40102
rect 116082 40046 116138 40102
rect 115958 39922 116014 39978
rect 116082 39922 116138 39978
rect 146678 40294 146734 40350
rect 146802 40294 146858 40350
rect 146678 40170 146734 40226
rect 146802 40170 146858 40226
rect 146678 40046 146734 40102
rect 146802 40046 146858 40102
rect 146678 39922 146734 39978
rect 146802 39922 146858 39978
rect 177398 40294 177454 40350
rect 177522 40294 177578 40350
rect 177398 40170 177454 40226
rect 177522 40170 177578 40226
rect 177398 40046 177454 40102
rect 177522 40046 177578 40102
rect 177398 39922 177454 39978
rect 177522 39922 177578 39978
rect 208118 40294 208174 40350
rect 208242 40294 208298 40350
rect 208118 40170 208174 40226
rect 208242 40170 208298 40226
rect 208118 40046 208174 40102
rect 208242 40046 208298 40102
rect 208118 39922 208174 39978
rect 208242 39922 208298 39978
rect 238838 40294 238894 40350
rect 238962 40294 239018 40350
rect 238838 40170 238894 40226
rect 238962 40170 239018 40226
rect 238838 40046 238894 40102
rect 238962 40046 239018 40102
rect 238838 39922 238894 39978
rect 238962 39922 239018 39978
rect 269558 40294 269614 40350
rect 269682 40294 269738 40350
rect 269558 40170 269614 40226
rect 269682 40170 269738 40226
rect 269558 40046 269614 40102
rect 269682 40046 269738 40102
rect 269558 39922 269614 39978
rect 269682 39922 269738 39978
rect 300278 40294 300334 40350
rect 300402 40294 300458 40350
rect 300278 40170 300334 40226
rect 300402 40170 300458 40226
rect 300278 40046 300334 40102
rect 300402 40046 300458 40102
rect 300278 39922 300334 39978
rect 300402 39922 300458 39978
rect 330998 40294 331054 40350
rect 331122 40294 331178 40350
rect 330998 40170 331054 40226
rect 331122 40170 331178 40226
rect 330998 40046 331054 40102
rect 331122 40046 331178 40102
rect 330998 39922 331054 39978
rect 331122 39922 331178 39978
rect 361718 40294 361774 40350
rect 361842 40294 361898 40350
rect 361718 40170 361774 40226
rect 361842 40170 361898 40226
rect 361718 40046 361774 40102
rect 361842 40046 361898 40102
rect 361718 39922 361774 39978
rect 361842 39922 361898 39978
rect 392438 40294 392494 40350
rect 392562 40294 392618 40350
rect 392438 40170 392494 40226
rect 392562 40170 392618 40226
rect 392438 40046 392494 40102
rect 392562 40046 392618 40102
rect 392438 39922 392494 39978
rect 392562 39922 392618 39978
rect 423158 40294 423214 40350
rect 423282 40294 423338 40350
rect 423158 40170 423214 40226
rect 423282 40170 423338 40226
rect 423158 40046 423214 40102
rect 423282 40046 423338 40102
rect 423158 39922 423214 39978
rect 423282 39922 423338 39978
rect 453878 40294 453934 40350
rect 454002 40294 454058 40350
rect 453878 40170 453934 40226
rect 454002 40170 454058 40226
rect 453878 40046 453934 40102
rect 454002 40046 454058 40102
rect 453878 39922 453934 39978
rect 454002 39922 454058 39978
rect 484598 40294 484654 40350
rect 484722 40294 484778 40350
rect 484598 40170 484654 40226
rect 484722 40170 484778 40226
rect 484598 40046 484654 40102
rect 484722 40046 484778 40102
rect 484598 39922 484654 39978
rect 484722 39922 484778 39978
rect 515318 40294 515374 40350
rect 515442 40294 515498 40350
rect 515318 40170 515374 40226
rect 515442 40170 515498 40226
rect 515318 40046 515374 40102
rect 515442 40046 515498 40102
rect 515318 39922 515374 39978
rect 515442 39922 515498 39978
rect 546038 40294 546094 40350
rect 546162 40294 546218 40350
rect 546038 40170 546094 40226
rect 546162 40170 546218 40226
rect 546038 40046 546094 40102
rect 546162 40046 546218 40102
rect 546038 39922 546094 39978
rect 546162 39922 546218 39978
rect 561250 40294 561306 40350
rect 561374 40294 561430 40350
rect 561498 40294 561554 40350
rect 561622 40294 561678 40350
rect 561250 40170 561306 40226
rect 561374 40170 561430 40226
rect 561498 40170 561554 40226
rect 561622 40170 561678 40226
rect 561250 40046 561306 40102
rect 561374 40046 561430 40102
rect 561498 40046 561554 40102
rect 561622 40046 561678 40102
rect 561250 39922 561306 39978
rect 561374 39922 561430 39978
rect 561498 39922 561554 39978
rect 561622 39922 561678 39978
rect 111250 22294 111306 22350
rect 111374 22294 111430 22350
rect 111498 22294 111554 22350
rect 111622 22294 111678 22350
rect 111250 22170 111306 22226
rect 111374 22170 111430 22226
rect 111498 22170 111554 22226
rect 111622 22170 111678 22226
rect 111250 22046 111306 22102
rect 111374 22046 111430 22102
rect 111498 22046 111554 22102
rect 111622 22046 111678 22102
rect 111250 21922 111306 21978
rect 111374 21922 111430 21978
rect 111498 21922 111554 21978
rect 111622 21922 111678 21978
rect 111250 4294 111306 4350
rect 111374 4294 111430 4350
rect 111498 4294 111554 4350
rect 111622 4294 111678 4350
rect 111250 4170 111306 4226
rect 111374 4170 111430 4226
rect 111498 4170 111554 4226
rect 111622 4170 111678 4226
rect 111250 4046 111306 4102
rect 111374 4046 111430 4102
rect 111498 4046 111554 4102
rect 111622 4046 111678 4102
rect 111250 3922 111306 3978
rect 111374 3922 111430 3978
rect 111498 3922 111554 3978
rect 111622 3922 111678 3978
rect 111250 -216 111306 -160
rect 111374 -216 111430 -160
rect 111498 -216 111554 -160
rect 111622 -216 111678 -160
rect 111250 -340 111306 -284
rect 111374 -340 111430 -284
rect 111498 -340 111554 -284
rect 111622 -340 111678 -284
rect 111250 -464 111306 -408
rect 111374 -464 111430 -408
rect 111498 -464 111554 -408
rect 111622 -464 111678 -408
rect 111250 -588 111306 -532
rect 111374 -588 111430 -532
rect 111498 -588 111554 -532
rect 111622 -588 111678 -532
rect 114970 28294 115026 28350
rect 115094 28294 115150 28350
rect 115218 28294 115274 28350
rect 115342 28294 115398 28350
rect 114970 28170 115026 28226
rect 115094 28170 115150 28226
rect 115218 28170 115274 28226
rect 115342 28170 115398 28226
rect 114970 28046 115026 28102
rect 115094 28046 115150 28102
rect 115218 28046 115274 28102
rect 115342 28046 115398 28102
rect 114970 27922 115026 27978
rect 115094 27922 115150 27978
rect 115218 27922 115274 27978
rect 115342 27922 115398 27978
rect 114970 10294 115026 10350
rect 115094 10294 115150 10350
rect 115218 10294 115274 10350
rect 115342 10294 115398 10350
rect 114970 10170 115026 10226
rect 115094 10170 115150 10226
rect 115218 10170 115274 10226
rect 115342 10170 115398 10226
rect 114970 10046 115026 10102
rect 115094 10046 115150 10102
rect 115218 10046 115274 10102
rect 115342 10046 115398 10102
rect 114970 9922 115026 9978
rect 115094 9922 115150 9978
rect 115218 9922 115274 9978
rect 115342 9922 115398 9978
rect 114970 -1176 115026 -1120
rect 115094 -1176 115150 -1120
rect 115218 -1176 115274 -1120
rect 115342 -1176 115398 -1120
rect 114970 -1300 115026 -1244
rect 115094 -1300 115150 -1244
rect 115218 -1300 115274 -1244
rect 115342 -1300 115398 -1244
rect 114970 -1424 115026 -1368
rect 115094 -1424 115150 -1368
rect 115218 -1424 115274 -1368
rect 115342 -1424 115398 -1368
rect 114970 -1548 115026 -1492
rect 115094 -1548 115150 -1492
rect 115218 -1548 115274 -1492
rect 115342 -1548 115398 -1492
rect 129250 22294 129306 22350
rect 129374 22294 129430 22350
rect 129498 22294 129554 22350
rect 129622 22294 129678 22350
rect 129250 22170 129306 22226
rect 129374 22170 129430 22226
rect 129498 22170 129554 22226
rect 129622 22170 129678 22226
rect 129250 22046 129306 22102
rect 129374 22046 129430 22102
rect 129498 22046 129554 22102
rect 129622 22046 129678 22102
rect 129250 21922 129306 21978
rect 129374 21922 129430 21978
rect 129498 21922 129554 21978
rect 129622 21922 129678 21978
rect 129250 4294 129306 4350
rect 129374 4294 129430 4350
rect 129498 4294 129554 4350
rect 129622 4294 129678 4350
rect 129250 4170 129306 4226
rect 129374 4170 129430 4226
rect 129498 4170 129554 4226
rect 129622 4170 129678 4226
rect 129250 4046 129306 4102
rect 129374 4046 129430 4102
rect 129498 4046 129554 4102
rect 129622 4046 129678 4102
rect 129250 3922 129306 3978
rect 129374 3922 129430 3978
rect 129498 3922 129554 3978
rect 129622 3922 129678 3978
rect 129250 -216 129306 -160
rect 129374 -216 129430 -160
rect 129498 -216 129554 -160
rect 129622 -216 129678 -160
rect 129250 -340 129306 -284
rect 129374 -340 129430 -284
rect 129498 -340 129554 -284
rect 129622 -340 129678 -284
rect 129250 -464 129306 -408
rect 129374 -464 129430 -408
rect 129498 -464 129554 -408
rect 129622 -464 129678 -408
rect 129250 -588 129306 -532
rect 129374 -588 129430 -532
rect 129498 -588 129554 -532
rect 129622 -588 129678 -532
rect 132970 28294 133026 28350
rect 133094 28294 133150 28350
rect 133218 28294 133274 28350
rect 133342 28294 133398 28350
rect 132970 28170 133026 28226
rect 133094 28170 133150 28226
rect 133218 28170 133274 28226
rect 133342 28170 133398 28226
rect 132970 28046 133026 28102
rect 133094 28046 133150 28102
rect 133218 28046 133274 28102
rect 133342 28046 133398 28102
rect 132970 27922 133026 27978
rect 133094 27922 133150 27978
rect 133218 27922 133274 27978
rect 133342 27922 133398 27978
rect 132970 10294 133026 10350
rect 133094 10294 133150 10350
rect 133218 10294 133274 10350
rect 133342 10294 133398 10350
rect 132970 10170 133026 10226
rect 133094 10170 133150 10226
rect 133218 10170 133274 10226
rect 133342 10170 133398 10226
rect 132970 10046 133026 10102
rect 133094 10046 133150 10102
rect 133218 10046 133274 10102
rect 133342 10046 133398 10102
rect 132970 9922 133026 9978
rect 133094 9922 133150 9978
rect 133218 9922 133274 9978
rect 133342 9922 133398 9978
rect 132970 -1176 133026 -1120
rect 133094 -1176 133150 -1120
rect 133218 -1176 133274 -1120
rect 133342 -1176 133398 -1120
rect 132970 -1300 133026 -1244
rect 133094 -1300 133150 -1244
rect 133218 -1300 133274 -1244
rect 133342 -1300 133398 -1244
rect 132970 -1424 133026 -1368
rect 133094 -1424 133150 -1368
rect 133218 -1424 133274 -1368
rect 133342 -1424 133398 -1368
rect 132970 -1548 133026 -1492
rect 133094 -1548 133150 -1492
rect 133218 -1548 133274 -1492
rect 133342 -1548 133398 -1492
rect 147250 22294 147306 22350
rect 147374 22294 147430 22350
rect 147498 22294 147554 22350
rect 147622 22294 147678 22350
rect 147250 22170 147306 22226
rect 147374 22170 147430 22226
rect 147498 22170 147554 22226
rect 147622 22170 147678 22226
rect 147250 22046 147306 22102
rect 147374 22046 147430 22102
rect 147498 22046 147554 22102
rect 147622 22046 147678 22102
rect 147250 21922 147306 21978
rect 147374 21922 147430 21978
rect 147498 21922 147554 21978
rect 147622 21922 147678 21978
rect 147250 4294 147306 4350
rect 147374 4294 147430 4350
rect 147498 4294 147554 4350
rect 147622 4294 147678 4350
rect 147250 4170 147306 4226
rect 147374 4170 147430 4226
rect 147498 4170 147554 4226
rect 147622 4170 147678 4226
rect 147250 4046 147306 4102
rect 147374 4046 147430 4102
rect 147498 4046 147554 4102
rect 147622 4046 147678 4102
rect 147250 3922 147306 3978
rect 147374 3922 147430 3978
rect 147498 3922 147554 3978
rect 147622 3922 147678 3978
rect 147250 -216 147306 -160
rect 147374 -216 147430 -160
rect 147498 -216 147554 -160
rect 147622 -216 147678 -160
rect 147250 -340 147306 -284
rect 147374 -340 147430 -284
rect 147498 -340 147554 -284
rect 147622 -340 147678 -284
rect 147250 -464 147306 -408
rect 147374 -464 147430 -408
rect 147498 -464 147554 -408
rect 147622 -464 147678 -408
rect 147250 -588 147306 -532
rect 147374 -588 147430 -532
rect 147498 -588 147554 -532
rect 147622 -588 147678 -532
rect 150970 28294 151026 28350
rect 151094 28294 151150 28350
rect 151218 28294 151274 28350
rect 151342 28294 151398 28350
rect 150970 28170 151026 28226
rect 151094 28170 151150 28226
rect 151218 28170 151274 28226
rect 151342 28170 151398 28226
rect 150970 28046 151026 28102
rect 151094 28046 151150 28102
rect 151218 28046 151274 28102
rect 151342 28046 151398 28102
rect 150970 27922 151026 27978
rect 151094 27922 151150 27978
rect 151218 27922 151274 27978
rect 151342 27922 151398 27978
rect 150970 10294 151026 10350
rect 151094 10294 151150 10350
rect 151218 10294 151274 10350
rect 151342 10294 151398 10350
rect 150970 10170 151026 10226
rect 151094 10170 151150 10226
rect 151218 10170 151274 10226
rect 151342 10170 151398 10226
rect 150970 10046 151026 10102
rect 151094 10046 151150 10102
rect 151218 10046 151274 10102
rect 151342 10046 151398 10102
rect 150970 9922 151026 9978
rect 151094 9922 151150 9978
rect 151218 9922 151274 9978
rect 151342 9922 151398 9978
rect 150970 -1176 151026 -1120
rect 151094 -1176 151150 -1120
rect 151218 -1176 151274 -1120
rect 151342 -1176 151398 -1120
rect 150970 -1300 151026 -1244
rect 151094 -1300 151150 -1244
rect 151218 -1300 151274 -1244
rect 151342 -1300 151398 -1244
rect 150970 -1424 151026 -1368
rect 151094 -1424 151150 -1368
rect 151218 -1424 151274 -1368
rect 151342 -1424 151398 -1368
rect 150970 -1548 151026 -1492
rect 151094 -1548 151150 -1492
rect 151218 -1548 151274 -1492
rect 151342 -1548 151398 -1492
rect 165250 22294 165306 22350
rect 165374 22294 165430 22350
rect 165498 22294 165554 22350
rect 165622 22294 165678 22350
rect 165250 22170 165306 22226
rect 165374 22170 165430 22226
rect 165498 22170 165554 22226
rect 165622 22170 165678 22226
rect 165250 22046 165306 22102
rect 165374 22046 165430 22102
rect 165498 22046 165554 22102
rect 165622 22046 165678 22102
rect 165250 21922 165306 21978
rect 165374 21922 165430 21978
rect 165498 21922 165554 21978
rect 165622 21922 165678 21978
rect 165250 4294 165306 4350
rect 165374 4294 165430 4350
rect 165498 4294 165554 4350
rect 165622 4294 165678 4350
rect 165250 4170 165306 4226
rect 165374 4170 165430 4226
rect 165498 4170 165554 4226
rect 165622 4170 165678 4226
rect 165250 4046 165306 4102
rect 165374 4046 165430 4102
rect 165498 4046 165554 4102
rect 165622 4046 165678 4102
rect 165250 3922 165306 3978
rect 165374 3922 165430 3978
rect 165498 3922 165554 3978
rect 165622 3922 165678 3978
rect 165250 -216 165306 -160
rect 165374 -216 165430 -160
rect 165498 -216 165554 -160
rect 165622 -216 165678 -160
rect 165250 -340 165306 -284
rect 165374 -340 165430 -284
rect 165498 -340 165554 -284
rect 165622 -340 165678 -284
rect 165250 -464 165306 -408
rect 165374 -464 165430 -408
rect 165498 -464 165554 -408
rect 165622 -464 165678 -408
rect 165250 -588 165306 -532
rect 165374 -588 165430 -532
rect 165498 -588 165554 -532
rect 165622 -588 165678 -532
rect 168970 28294 169026 28350
rect 169094 28294 169150 28350
rect 169218 28294 169274 28350
rect 169342 28294 169398 28350
rect 168970 28170 169026 28226
rect 169094 28170 169150 28226
rect 169218 28170 169274 28226
rect 169342 28170 169398 28226
rect 168970 28046 169026 28102
rect 169094 28046 169150 28102
rect 169218 28046 169274 28102
rect 169342 28046 169398 28102
rect 168970 27922 169026 27978
rect 169094 27922 169150 27978
rect 169218 27922 169274 27978
rect 169342 27922 169398 27978
rect 168970 10294 169026 10350
rect 169094 10294 169150 10350
rect 169218 10294 169274 10350
rect 169342 10294 169398 10350
rect 168970 10170 169026 10226
rect 169094 10170 169150 10226
rect 169218 10170 169274 10226
rect 169342 10170 169398 10226
rect 168970 10046 169026 10102
rect 169094 10046 169150 10102
rect 169218 10046 169274 10102
rect 169342 10046 169398 10102
rect 168970 9922 169026 9978
rect 169094 9922 169150 9978
rect 169218 9922 169274 9978
rect 169342 9922 169398 9978
rect 168970 -1176 169026 -1120
rect 169094 -1176 169150 -1120
rect 169218 -1176 169274 -1120
rect 169342 -1176 169398 -1120
rect 168970 -1300 169026 -1244
rect 169094 -1300 169150 -1244
rect 169218 -1300 169274 -1244
rect 169342 -1300 169398 -1244
rect 168970 -1424 169026 -1368
rect 169094 -1424 169150 -1368
rect 169218 -1424 169274 -1368
rect 169342 -1424 169398 -1368
rect 168970 -1548 169026 -1492
rect 169094 -1548 169150 -1492
rect 169218 -1548 169274 -1492
rect 169342 -1548 169398 -1492
rect 183250 22294 183306 22350
rect 183374 22294 183430 22350
rect 183498 22294 183554 22350
rect 183622 22294 183678 22350
rect 183250 22170 183306 22226
rect 183374 22170 183430 22226
rect 183498 22170 183554 22226
rect 183622 22170 183678 22226
rect 183250 22046 183306 22102
rect 183374 22046 183430 22102
rect 183498 22046 183554 22102
rect 183622 22046 183678 22102
rect 183250 21922 183306 21978
rect 183374 21922 183430 21978
rect 183498 21922 183554 21978
rect 183622 21922 183678 21978
rect 183250 4294 183306 4350
rect 183374 4294 183430 4350
rect 183498 4294 183554 4350
rect 183622 4294 183678 4350
rect 183250 4170 183306 4226
rect 183374 4170 183430 4226
rect 183498 4170 183554 4226
rect 183622 4170 183678 4226
rect 183250 4046 183306 4102
rect 183374 4046 183430 4102
rect 183498 4046 183554 4102
rect 183622 4046 183678 4102
rect 183250 3922 183306 3978
rect 183374 3922 183430 3978
rect 183498 3922 183554 3978
rect 183622 3922 183678 3978
rect 183250 -216 183306 -160
rect 183374 -216 183430 -160
rect 183498 -216 183554 -160
rect 183622 -216 183678 -160
rect 183250 -340 183306 -284
rect 183374 -340 183430 -284
rect 183498 -340 183554 -284
rect 183622 -340 183678 -284
rect 183250 -464 183306 -408
rect 183374 -464 183430 -408
rect 183498 -464 183554 -408
rect 183622 -464 183678 -408
rect 183250 -588 183306 -532
rect 183374 -588 183430 -532
rect 183498 -588 183554 -532
rect 183622 -588 183678 -532
rect 186970 28294 187026 28350
rect 187094 28294 187150 28350
rect 187218 28294 187274 28350
rect 187342 28294 187398 28350
rect 186970 28170 187026 28226
rect 187094 28170 187150 28226
rect 187218 28170 187274 28226
rect 187342 28170 187398 28226
rect 186970 28046 187026 28102
rect 187094 28046 187150 28102
rect 187218 28046 187274 28102
rect 187342 28046 187398 28102
rect 186970 27922 187026 27978
rect 187094 27922 187150 27978
rect 187218 27922 187274 27978
rect 187342 27922 187398 27978
rect 186970 10294 187026 10350
rect 187094 10294 187150 10350
rect 187218 10294 187274 10350
rect 187342 10294 187398 10350
rect 186970 10170 187026 10226
rect 187094 10170 187150 10226
rect 187218 10170 187274 10226
rect 187342 10170 187398 10226
rect 186970 10046 187026 10102
rect 187094 10046 187150 10102
rect 187218 10046 187274 10102
rect 187342 10046 187398 10102
rect 186970 9922 187026 9978
rect 187094 9922 187150 9978
rect 187218 9922 187274 9978
rect 187342 9922 187398 9978
rect 186970 -1176 187026 -1120
rect 187094 -1176 187150 -1120
rect 187218 -1176 187274 -1120
rect 187342 -1176 187398 -1120
rect 186970 -1300 187026 -1244
rect 187094 -1300 187150 -1244
rect 187218 -1300 187274 -1244
rect 187342 -1300 187398 -1244
rect 186970 -1424 187026 -1368
rect 187094 -1424 187150 -1368
rect 187218 -1424 187274 -1368
rect 187342 -1424 187398 -1368
rect 186970 -1548 187026 -1492
rect 187094 -1548 187150 -1492
rect 187218 -1548 187274 -1492
rect 187342 -1548 187398 -1492
rect 201250 22294 201306 22350
rect 201374 22294 201430 22350
rect 201498 22294 201554 22350
rect 201622 22294 201678 22350
rect 201250 22170 201306 22226
rect 201374 22170 201430 22226
rect 201498 22170 201554 22226
rect 201622 22170 201678 22226
rect 201250 22046 201306 22102
rect 201374 22046 201430 22102
rect 201498 22046 201554 22102
rect 201622 22046 201678 22102
rect 201250 21922 201306 21978
rect 201374 21922 201430 21978
rect 201498 21922 201554 21978
rect 201622 21922 201678 21978
rect 201250 4294 201306 4350
rect 201374 4294 201430 4350
rect 201498 4294 201554 4350
rect 201622 4294 201678 4350
rect 201250 4170 201306 4226
rect 201374 4170 201430 4226
rect 201498 4170 201554 4226
rect 201622 4170 201678 4226
rect 201250 4046 201306 4102
rect 201374 4046 201430 4102
rect 201498 4046 201554 4102
rect 201622 4046 201678 4102
rect 201250 3922 201306 3978
rect 201374 3922 201430 3978
rect 201498 3922 201554 3978
rect 201622 3922 201678 3978
rect 201250 -216 201306 -160
rect 201374 -216 201430 -160
rect 201498 -216 201554 -160
rect 201622 -216 201678 -160
rect 201250 -340 201306 -284
rect 201374 -340 201430 -284
rect 201498 -340 201554 -284
rect 201622 -340 201678 -284
rect 201250 -464 201306 -408
rect 201374 -464 201430 -408
rect 201498 -464 201554 -408
rect 201622 -464 201678 -408
rect 201250 -588 201306 -532
rect 201374 -588 201430 -532
rect 201498 -588 201554 -532
rect 201622 -588 201678 -532
rect 204970 28294 205026 28350
rect 205094 28294 205150 28350
rect 205218 28294 205274 28350
rect 205342 28294 205398 28350
rect 204970 28170 205026 28226
rect 205094 28170 205150 28226
rect 205218 28170 205274 28226
rect 205342 28170 205398 28226
rect 204970 28046 205026 28102
rect 205094 28046 205150 28102
rect 205218 28046 205274 28102
rect 205342 28046 205398 28102
rect 204970 27922 205026 27978
rect 205094 27922 205150 27978
rect 205218 27922 205274 27978
rect 205342 27922 205398 27978
rect 204970 10294 205026 10350
rect 205094 10294 205150 10350
rect 205218 10294 205274 10350
rect 205342 10294 205398 10350
rect 204970 10170 205026 10226
rect 205094 10170 205150 10226
rect 205218 10170 205274 10226
rect 205342 10170 205398 10226
rect 204970 10046 205026 10102
rect 205094 10046 205150 10102
rect 205218 10046 205274 10102
rect 205342 10046 205398 10102
rect 204970 9922 205026 9978
rect 205094 9922 205150 9978
rect 205218 9922 205274 9978
rect 205342 9922 205398 9978
rect 204970 -1176 205026 -1120
rect 205094 -1176 205150 -1120
rect 205218 -1176 205274 -1120
rect 205342 -1176 205398 -1120
rect 204970 -1300 205026 -1244
rect 205094 -1300 205150 -1244
rect 205218 -1300 205274 -1244
rect 205342 -1300 205398 -1244
rect 204970 -1424 205026 -1368
rect 205094 -1424 205150 -1368
rect 205218 -1424 205274 -1368
rect 205342 -1424 205398 -1368
rect 204970 -1548 205026 -1492
rect 205094 -1548 205150 -1492
rect 205218 -1548 205274 -1492
rect 205342 -1548 205398 -1492
rect 219250 22294 219306 22350
rect 219374 22294 219430 22350
rect 219498 22294 219554 22350
rect 219622 22294 219678 22350
rect 219250 22170 219306 22226
rect 219374 22170 219430 22226
rect 219498 22170 219554 22226
rect 219622 22170 219678 22226
rect 219250 22046 219306 22102
rect 219374 22046 219430 22102
rect 219498 22046 219554 22102
rect 219622 22046 219678 22102
rect 219250 21922 219306 21978
rect 219374 21922 219430 21978
rect 219498 21922 219554 21978
rect 219622 21922 219678 21978
rect 219250 4294 219306 4350
rect 219374 4294 219430 4350
rect 219498 4294 219554 4350
rect 219622 4294 219678 4350
rect 219250 4170 219306 4226
rect 219374 4170 219430 4226
rect 219498 4170 219554 4226
rect 219622 4170 219678 4226
rect 219250 4046 219306 4102
rect 219374 4046 219430 4102
rect 219498 4046 219554 4102
rect 219622 4046 219678 4102
rect 219250 3922 219306 3978
rect 219374 3922 219430 3978
rect 219498 3922 219554 3978
rect 219622 3922 219678 3978
rect 219250 -216 219306 -160
rect 219374 -216 219430 -160
rect 219498 -216 219554 -160
rect 219622 -216 219678 -160
rect 219250 -340 219306 -284
rect 219374 -340 219430 -284
rect 219498 -340 219554 -284
rect 219622 -340 219678 -284
rect 219250 -464 219306 -408
rect 219374 -464 219430 -408
rect 219498 -464 219554 -408
rect 219622 -464 219678 -408
rect 219250 -588 219306 -532
rect 219374 -588 219430 -532
rect 219498 -588 219554 -532
rect 219622 -588 219678 -532
rect 222970 28294 223026 28350
rect 223094 28294 223150 28350
rect 223218 28294 223274 28350
rect 223342 28294 223398 28350
rect 222970 28170 223026 28226
rect 223094 28170 223150 28226
rect 223218 28170 223274 28226
rect 223342 28170 223398 28226
rect 222970 28046 223026 28102
rect 223094 28046 223150 28102
rect 223218 28046 223274 28102
rect 223342 28046 223398 28102
rect 222970 27922 223026 27978
rect 223094 27922 223150 27978
rect 223218 27922 223274 27978
rect 223342 27922 223398 27978
rect 222970 10294 223026 10350
rect 223094 10294 223150 10350
rect 223218 10294 223274 10350
rect 223342 10294 223398 10350
rect 222970 10170 223026 10226
rect 223094 10170 223150 10226
rect 223218 10170 223274 10226
rect 223342 10170 223398 10226
rect 222970 10046 223026 10102
rect 223094 10046 223150 10102
rect 223218 10046 223274 10102
rect 223342 10046 223398 10102
rect 222970 9922 223026 9978
rect 223094 9922 223150 9978
rect 223218 9922 223274 9978
rect 223342 9922 223398 9978
rect 222970 -1176 223026 -1120
rect 223094 -1176 223150 -1120
rect 223218 -1176 223274 -1120
rect 223342 -1176 223398 -1120
rect 222970 -1300 223026 -1244
rect 223094 -1300 223150 -1244
rect 223218 -1300 223274 -1244
rect 223342 -1300 223398 -1244
rect 222970 -1424 223026 -1368
rect 223094 -1424 223150 -1368
rect 223218 -1424 223274 -1368
rect 223342 -1424 223398 -1368
rect 222970 -1548 223026 -1492
rect 223094 -1548 223150 -1492
rect 223218 -1548 223274 -1492
rect 223342 -1548 223398 -1492
rect 237250 22294 237306 22350
rect 237374 22294 237430 22350
rect 237498 22294 237554 22350
rect 237622 22294 237678 22350
rect 237250 22170 237306 22226
rect 237374 22170 237430 22226
rect 237498 22170 237554 22226
rect 237622 22170 237678 22226
rect 237250 22046 237306 22102
rect 237374 22046 237430 22102
rect 237498 22046 237554 22102
rect 237622 22046 237678 22102
rect 237250 21922 237306 21978
rect 237374 21922 237430 21978
rect 237498 21922 237554 21978
rect 237622 21922 237678 21978
rect 237250 4294 237306 4350
rect 237374 4294 237430 4350
rect 237498 4294 237554 4350
rect 237622 4294 237678 4350
rect 237250 4170 237306 4226
rect 237374 4170 237430 4226
rect 237498 4170 237554 4226
rect 237622 4170 237678 4226
rect 237250 4046 237306 4102
rect 237374 4046 237430 4102
rect 237498 4046 237554 4102
rect 237622 4046 237678 4102
rect 237250 3922 237306 3978
rect 237374 3922 237430 3978
rect 237498 3922 237554 3978
rect 237622 3922 237678 3978
rect 237250 -216 237306 -160
rect 237374 -216 237430 -160
rect 237498 -216 237554 -160
rect 237622 -216 237678 -160
rect 237250 -340 237306 -284
rect 237374 -340 237430 -284
rect 237498 -340 237554 -284
rect 237622 -340 237678 -284
rect 237250 -464 237306 -408
rect 237374 -464 237430 -408
rect 237498 -464 237554 -408
rect 237622 -464 237678 -408
rect 237250 -588 237306 -532
rect 237374 -588 237430 -532
rect 237498 -588 237554 -532
rect 237622 -588 237678 -532
rect 240970 28294 241026 28350
rect 241094 28294 241150 28350
rect 241218 28294 241274 28350
rect 241342 28294 241398 28350
rect 240970 28170 241026 28226
rect 241094 28170 241150 28226
rect 241218 28170 241274 28226
rect 241342 28170 241398 28226
rect 240970 28046 241026 28102
rect 241094 28046 241150 28102
rect 241218 28046 241274 28102
rect 241342 28046 241398 28102
rect 240970 27922 241026 27978
rect 241094 27922 241150 27978
rect 241218 27922 241274 27978
rect 241342 27922 241398 27978
rect 240970 10294 241026 10350
rect 241094 10294 241150 10350
rect 241218 10294 241274 10350
rect 241342 10294 241398 10350
rect 240970 10170 241026 10226
rect 241094 10170 241150 10226
rect 241218 10170 241274 10226
rect 241342 10170 241398 10226
rect 240970 10046 241026 10102
rect 241094 10046 241150 10102
rect 241218 10046 241274 10102
rect 241342 10046 241398 10102
rect 240970 9922 241026 9978
rect 241094 9922 241150 9978
rect 241218 9922 241274 9978
rect 241342 9922 241398 9978
rect 240970 -1176 241026 -1120
rect 241094 -1176 241150 -1120
rect 241218 -1176 241274 -1120
rect 241342 -1176 241398 -1120
rect 240970 -1300 241026 -1244
rect 241094 -1300 241150 -1244
rect 241218 -1300 241274 -1244
rect 241342 -1300 241398 -1244
rect 240970 -1424 241026 -1368
rect 241094 -1424 241150 -1368
rect 241218 -1424 241274 -1368
rect 241342 -1424 241398 -1368
rect 240970 -1548 241026 -1492
rect 241094 -1548 241150 -1492
rect 241218 -1548 241274 -1492
rect 241342 -1548 241398 -1492
rect 255250 22294 255306 22350
rect 255374 22294 255430 22350
rect 255498 22294 255554 22350
rect 255622 22294 255678 22350
rect 255250 22170 255306 22226
rect 255374 22170 255430 22226
rect 255498 22170 255554 22226
rect 255622 22170 255678 22226
rect 255250 22046 255306 22102
rect 255374 22046 255430 22102
rect 255498 22046 255554 22102
rect 255622 22046 255678 22102
rect 255250 21922 255306 21978
rect 255374 21922 255430 21978
rect 255498 21922 255554 21978
rect 255622 21922 255678 21978
rect 255250 4294 255306 4350
rect 255374 4294 255430 4350
rect 255498 4294 255554 4350
rect 255622 4294 255678 4350
rect 255250 4170 255306 4226
rect 255374 4170 255430 4226
rect 255498 4170 255554 4226
rect 255622 4170 255678 4226
rect 255250 4046 255306 4102
rect 255374 4046 255430 4102
rect 255498 4046 255554 4102
rect 255622 4046 255678 4102
rect 255250 3922 255306 3978
rect 255374 3922 255430 3978
rect 255498 3922 255554 3978
rect 255622 3922 255678 3978
rect 255250 -216 255306 -160
rect 255374 -216 255430 -160
rect 255498 -216 255554 -160
rect 255622 -216 255678 -160
rect 255250 -340 255306 -284
rect 255374 -340 255430 -284
rect 255498 -340 255554 -284
rect 255622 -340 255678 -284
rect 255250 -464 255306 -408
rect 255374 -464 255430 -408
rect 255498 -464 255554 -408
rect 255622 -464 255678 -408
rect 255250 -588 255306 -532
rect 255374 -588 255430 -532
rect 255498 -588 255554 -532
rect 255622 -588 255678 -532
rect 258970 28294 259026 28350
rect 259094 28294 259150 28350
rect 259218 28294 259274 28350
rect 259342 28294 259398 28350
rect 258970 28170 259026 28226
rect 259094 28170 259150 28226
rect 259218 28170 259274 28226
rect 259342 28170 259398 28226
rect 258970 28046 259026 28102
rect 259094 28046 259150 28102
rect 259218 28046 259274 28102
rect 259342 28046 259398 28102
rect 258970 27922 259026 27978
rect 259094 27922 259150 27978
rect 259218 27922 259274 27978
rect 259342 27922 259398 27978
rect 258970 10294 259026 10350
rect 259094 10294 259150 10350
rect 259218 10294 259274 10350
rect 259342 10294 259398 10350
rect 258970 10170 259026 10226
rect 259094 10170 259150 10226
rect 259218 10170 259274 10226
rect 259342 10170 259398 10226
rect 258970 10046 259026 10102
rect 259094 10046 259150 10102
rect 259218 10046 259274 10102
rect 259342 10046 259398 10102
rect 258970 9922 259026 9978
rect 259094 9922 259150 9978
rect 259218 9922 259274 9978
rect 259342 9922 259398 9978
rect 258970 -1176 259026 -1120
rect 259094 -1176 259150 -1120
rect 259218 -1176 259274 -1120
rect 259342 -1176 259398 -1120
rect 258970 -1300 259026 -1244
rect 259094 -1300 259150 -1244
rect 259218 -1300 259274 -1244
rect 259342 -1300 259398 -1244
rect 258970 -1424 259026 -1368
rect 259094 -1424 259150 -1368
rect 259218 -1424 259274 -1368
rect 259342 -1424 259398 -1368
rect 258970 -1548 259026 -1492
rect 259094 -1548 259150 -1492
rect 259218 -1548 259274 -1492
rect 259342 -1548 259398 -1492
rect 273250 22294 273306 22350
rect 273374 22294 273430 22350
rect 273498 22294 273554 22350
rect 273622 22294 273678 22350
rect 273250 22170 273306 22226
rect 273374 22170 273430 22226
rect 273498 22170 273554 22226
rect 273622 22170 273678 22226
rect 273250 22046 273306 22102
rect 273374 22046 273430 22102
rect 273498 22046 273554 22102
rect 273622 22046 273678 22102
rect 273250 21922 273306 21978
rect 273374 21922 273430 21978
rect 273498 21922 273554 21978
rect 273622 21922 273678 21978
rect 273250 4294 273306 4350
rect 273374 4294 273430 4350
rect 273498 4294 273554 4350
rect 273622 4294 273678 4350
rect 273250 4170 273306 4226
rect 273374 4170 273430 4226
rect 273498 4170 273554 4226
rect 273622 4170 273678 4226
rect 273250 4046 273306 4102
rect 273374 4046 273430 4102
rect 273498 4046 273554 4102
rect 273622 4046 273678 4102
rect 273250 3922 273306 3978
rect 273374 3922 273430 3978
rect 273498 3922 273554 3978
rect 273622 3922 273678 3978
rect 273250 -216 273306 -160
rect 273374 -216 273430 -160
rect 273498 -216 273554 -160
rect 273622 -216 273678 -160
rect 273250 -340 273306 -284
rect 273374 -340 273430 -284
rect 273498 -340 273554 -284
rect 273622 -340 273678 -284
rect 273250 -464 273306 -408
rect 273374 -464 273430 -408
rect 273498 -464 273554 -408
rect 273622 -464 273678 -408
rect 273250 -588 273306 -532
rect 273374 -588 273430 -532
rect 273498 -588 273554 -532
rect 273622 -588 273678 -532
rect 276970 28294 277026 28350
rect 277094 28294 277150 28350
rect 277218 28294 277274 28350
rect 277342 28294 277398 28350
rect 276970 28170 277026 28226
rect 277094 28170 277150 28226
rect 277218 28170 277274 28226
rect 277342 28170 277398 28226
rect 276970 28046 277026 28102
rect 277094 28046 277150 28102
rect 277218 28046 277274 28102
rect 277342 28046 277398 28102
rect 276970 27922 277026 27978
rect 277094 27922 277150 27978
rect 277218 27922 277274 27978
rect 277342 27922 277398 27978
rect 276970 10294 277026 10350
rect 277094 10294 277150 10350
rect 277218 10294 277274 10350
rect 277342 10294 277398 10350
rect 276970 10170 277026 10226
rect 277094 10170 277150 10226
rect 277218 10170 277274 10226
rect 277342 10170 277398 10226
rect 276970 10046 277026 10102
rect 277094 10046 277150 10102
rect 277218 10046 277274 10102
rect 277342 10046 277398 10102
rect 276970 9922 277026 9978
rect 277094 9922 277150 9978
rect 277218 9922 277274 9978
rect 277342 9922 277398 9978
rect 276970 -1176 277026 -1120
rect 277094 -1176 277150 -1120
rect 277218 -1176 277274 -1120
rect 277342 -1176 277398 -1120
rect 276970 -1300 277026 -1244
rect 277094 -1300 277150 -1244
rect 277218 -1300 277274 -1244
rect 277342 -1300 277398 -1244
rect 276970 -1424 277026 -1368
rect 277094 -1424 277150 -1368
rect 277218 -1424 277274 -1368
rect 277342 -1424 277398 -1368
rect 276970 -1548 277026 -1492
rect 277094 -1548 277150 -1492
rect 277218 -1548 277274 -1492
rect 277342 -1548 277398 -1492
rect 291250 22294 291306 22350
rect 291374 22294 291430 22350
rect 291498 22294 291554 22350
rect 291622 22294 291678 22350
rect 291250 22170 291306 22226
rect 291374 22170 291430 22226
rect 291498 22170 291554 22226
rect 291622 22170 291678 22226
rect 291250 22046 291306 22102
rect 291374 22046 291430 22102
rect 291498 22046 291554 22102
rect 291622 22046 291678 22102
rect 291250 21922 291306 21978
rect 291374 21922 291430 21978
rect 291498 21922 291554 21978
rect 291622 21922 291678 21978
rect 291250 4294 291306 4350
rect 291374 4294 291430 4350
rect 291498 4294 291554 4350
rect 291622 4294 291678 4350
rect 291250 4170 291306 4226
rect 291374 4170 291430 4226
rect 291498 4170 291554 4226
rect 291622 4170 291678 4226
rect 291250 4046 291306 4102
rect 291374 4046 291430 4102
rect 291498 4046 291554 4102
rect 291622 4046 291678 4102
rect 291250 3922 291306 3978
rect 291374 3922 291430 3978
rect 291498 3922 291554 3978
rect 291622 3922 291678 3978
rect 291250 -216 291306 -160
rect 291374 -216 291430 -160
rect 291498 -216 291554 -160
rect 291622 -216 291678 -160
rect 291250 -340 291306 -284
rect 291374 -340 291430 -284
rect 291498 -340 291554 -284
rect 291622 -340 291678 -284
rect 291250 -464 291306 -408
rect 291374 -464 291430 -408
rect 291498 -464 291554 -408
rect 291622 -464 291678 -408
rect 291250 -588 291306 -532
rect 291374 -588 291430 -532
rect 291498 -588 291554 -532
rect 291622 -588 291678 -532
rect 294970 28294 295026 28350
rect 295094 28294 295150 28350
rect 295218 28294 295274 28350
rect 295342 28294 295398 28350
rect 294970 28170 295026 28226
rect 295094 28170 295150 28226
rect 295218 28170 295274 28226
rect 295342 28170 295398 28226
rect 294970 28046 295026 28102
rect 295094 28046 295150 28102
rect 295218 28046 295274 28102
rect 295342 28046 295398 28102
rect 294970 27922 295026 27978
rect 295094 27922 295150 27978
rect 295218 27922 295274 27978
rect 295342 27922 295398 27978
rect 294970 10294 295026 10350
rect 295094 10294 295150 10350
rect 295218 10294 295274 10350
rect 295342 10294 295398 10350
rect 294970 10170 295026 10226
rect 295094 10170 295150 10226
rect 295218 10170 295274 10226
rect 295342 10170 295398 10226
rect 294970 10046 295026 10102
rect 295094 10046 295150 10102
rect 295218 10046 295274 10102
rect 295342 10046 295398 10102
rect 294970 9922 295026 9978
rect 295094 9922 295150 9978
rect 295218 9922 295274 9978
rect 295342 9922 295398 9978
rect 294970 -1176 295026 -1120
rect 295094 -1176 295150 -1120
rect 295218 -1176 295274 -1120
rect 295342 -1176 295398 -1120
rect 294970 -1300 295026 -1244
rect 295094 -1300 295150 -1244
rect 295218 -1300 295274 -1244
rect 295342 -1300 295398 -1244
rect 294970 -1424 295026 -1368
rect 295094 -1424 295150 -1368
rect 295218 -1424 295274 -1368
rect 295342 -1424 295398 -1368
rect 294970 -1548 295026 -1492
rect 295094 -1548 295150 -1492
rect 295218 -1548 295274 -1492
rect 295342 -1548 295398 -1492
rect 309250 22294 309306 22350
rect 309374 22294 309430 22350
rect 309498 22294 309554 22350
rect 309622 22294 309678 22350
rect 309250 22170 309306 22226
rect 309374 22170 309430 22226
rect 309498 22170 309554 22226
rect 309622 22170 309678 22226
rect 309250 22046 309306 22102
rect 309374 22046 309430 22102
rect 309498 22046 309554 22102
rect 309622 22046 309678 22102
rect 309250 21922 309306 21978
rect 309374 21922 309430 21978
rect 309498 21922 309554 21978
rect 309622 21922 309678 21978
rect 309250 4294 309306 4350
rect 309374 4294 309430 4350
rect 309498 4294 309554 4350
rect 309622 4294 309678 4350
rect 309250 4170 309306 4226
rect 309374 4170 309430 4226
rect 309498 4170 309554 4226
rect 309622 4170 309678 4226
rect 309250 4046 309306 4102
rect 309374 4046 309430 4102
rect 309498 4046 309554 4102
rect 309622 4046 309678 4102
rect 309250 3922 309306 3978
rect 309374 3922 309430 3978
rect 309498 3922 309554 3978
rect 309622 3922 309678 3978
rect 309250 -216 309306 -160
rect 309374 -216 309430 -160
rect 309498 -216 309554 -160
rect 309622 -216 309678 -160
rect 309250 -340 309306 -284
rect 309374 -340 309430 -284
rect 309498 -340 309554 -284
rect 309622 -340 309678 -284
rect 309250 -464 309306 -408
rect 309374 -464 309430 -408
rect 309498 -464 309554 -408
rect 309622 -464 309678 -408
rect 309250 -588 309306 -532
rect 309374 -588 309430 -532
rect 309498 -588 309554 -532
rect 309622 -588 309678 -532
rect 312970 28294 313026 28350
rect 313094 28294 313150 28350
rect 313218 28294 313274 28350
rect 313342 28294 313398 28350
rect 312970 28170 313026 28226
rect 313094 28170 313150 28226
rect 313218 28170 313274 28226
rect 313342 28170 313398 28226
rect 312970 28046 313026 28102
rect 313094 28046 313150 28102
rect 313218 28046 313274 28102
rect 313342 28046 313398 28102
rect 312970 27922 313026 27978
rect 313094 27922 313150 27978
rect 313218 27922 313274 27978
rect 313342 27922 313398 27978
rect 312970 10294 313026 10350
rect 313094 10294 313150 10350
rect 313218 10294 313274 10350
rect 313342 10294 313398 10350
rect 312970 10170 313026 10226
rect 313094 10170 313150 10226
rect 313218 10170 313274 10226
rect 313342 10170 313398 10226
rect 312970 10046 313026 10102
rect 313094 10046 313150 10102
rect 313218 10046 313274 10102
rect 313342 10046 313398 10102
rect 312970 9922 313026 9978
rect 313094 9922 313150 9978
rect 313218 9922 313274 9978
rect 313342 9922 313398 9978
rect 312970 -1176 313026 -1120
rect 313094 -1176 313150 -1120
rect 313218 -1176 313274 -1120
rect 313342 -1176 313398 -1120
rect 312970 -1300 313026 -1244
rect 313094 -1300 313150 -1244
rect 313218 -1300 313274 -1244
rect 313342 -1300 313398 -1244
rect 312970 -1424 313026 -1368
rect 313094 -1424 313150 -1368
rect 313218 -1424 313274 -1368
rect 313342 -1424 313398 -1368
rect 312970 -1548 313026 -1492
rect 313094 -1548 313150 -1492
rect 313218 -1548 313274 -1492
rect 313342 -1548 313398 -1492
rect 327250 22294 327306 22350
rect 327374 22294 327430 22350
rect 327498 22294 327554 22350
rect 327622 22294 327678 22350
rect 327250 22170 327306 22226
rect 327374 22170 327430 22226
rect 327498 22170 327554 22226
rect 327622 22170 327678 22226
rect 327250 22046 327306 22102
rect 327374 22046 327430 22102
rect 327498 22046 327554 22102
rect 327622 22046 327678 22102
rect 327250 21922 327306 21978
rect 327374 21922 327430 21978
rect 327498 21922 327554 21978
rect 327622 21922 327678 21978
rect 327250 4294 327306 4350
rect 327374 4294 327430 4350
rect 327498 4294 327554 4350
rect 327622 4294 327678 4350
rect 327250 4170 327306 4226
rect 327374 4170 327430 4226
rect 327498 4170 327554 4226
rect 327622 4170 327678 4226
rect 327250 4046 327306 4102
rect 327374 4046 327430 4102
rect 327498 4046 327554 4102
rect 327622 4046 327678 4102
rect 327250 3922 327306 3978
rect 327374 3922 327430 3978
rect 327498 3922 327554 3978
rect 327622 3922 327678 3978
rect 327250 -216 327306 -160
rect 327374 -216 327430 -160
rect 327498 -216 327554 -160
rect 327622 -216 327678 -160
rect 327250 -340 327306 -284
rect 327374 -340 327430 -284
rect 327498 -340 327554 -284
rect 327622 -340 327678 -284
rect 327250 -464 327306 -408
rect 327374 -464 327430 -408
rect 327498 -464 327554 -408
rect 327622 -464 327678 -408
rect 327250 -588 327306 -532
rect 327374 -588 327430 -532
rect 327498 -588 327554 -532
rect 327622 -588 327678 -532
rect 330970 28294 331026 28350
rect 331094 28294 331150 28350
rect 331218 28294 331274 28350
rect 331342 28294 331398 28350
rect 330970 28170 331026 28226
rect 331094 28170 331150 28226
rect 331218 28170 331274 28226
rect 331342 28170 331398 28226
rect 330970 28046 331026 28102
rect 331094 28046 331150 28102
rect 331218 28046 331274 28102
rect 331342 28046 331398 28102
rect 330970 27922 331026 27978
rect 331094 27922 331150 27978
rect 331218 27922 331274 27978
rect 331342 27922 331398 27978
rect 330970 10294 331026 10350
rect 331094 10294 331150 10350
rect 331218 10294 331274 10350
rect 331342 10294 331398 10350
rect 330970 10170 331026 10226
rect 331094 10170 331150 10226
rect 331218 10170 331274 10226
rect 331342 10170 331398 10226
rect 330970 10046 331026 10102
rect 331094 10046 331150 10102
rect 331218 10046 331274 10102
rect 331342 10046 331398 10102
rect 330970 9922 331026 9978
rect 331094 9922 331150 9978
rect 331218 9922 331274 9978
rect 331342 9922 331398 9978
rect 330970 -1176 331026 -1120
rect 331094 -1176 331150 -1120
rect 331218 -1176 331274 -1120
rect 331342 -1176 331398 -1120
rect 330970 -1300 331026 -1244
rect 331094 -1300 331150 -1244
rect 331218 -1300 331274 -1244
rect 331342 -1300 331398 -1244
rect 330970 -1424 331026 -1368
rect 331094 -1424 331150 -1368
rect 331218 -1424 331274 -1368
rect 331342 -1424 331398 -1368
rect 330970 -1548 331026 -1492
rect 331094 -1548 331150 -1492
rect 331218 -1548 331274 -1492
rect 331342 -1548 331398 -1492
rect 345250 22294 345306 22350
rect 345374 22294 345430 22350
rect 345498 22294 345554 22350
rect 345622 22294 345678 22350
rect 345250 22170 345306 22226
rect 345374 22170 345430 22226
rect 345498 22170 345554 22226
rect 345622 22170 345678 22226
rect 345250 22046 345306 22102
rect 345374 22046 345430 22102
rect 345498 22046 345554 22102
rect 345622 22046 345678 22102
rect 345250 21922 345306 21978
rect 345374 21922 345430 21978
rect 345498 21922 345554 21978
rect 345622 21922 345678 21978
rect 345250 4294 345306 4350
rect 345374 4294 345430 4350
rect 345498 4294 345554 4350
rect 345622 4294 345678 4350
rect 345250 4170 345306 4226
rect 345374 4170 345430 4226
rect 345498 4170 345554 4226
rect 345622 4170 345678 4226
rect 345250 4046 345306 4102
rect 345374 4046 345430 4102
rect 345498 4046 345554 4102
rect 345622 4046 345678 4102
rect 345250 3922 345306 3978
rect 345374 3922 345430 3978
rect 345498 3922 345554 3978
rect 345622 3922 345678 3978
rect 345250 -216 345306 -160
rect 345374 -216 345430 -160
rect 345498 -216 345554 -160
rect 345622 -216 345678 -160
rect 345250 -340 345306 -284
rect 345374 -340 345430 -284
rect 345498 -340 345554 -284
rect 345622 -340 345678 -284
rect 345250 -464 345306 -408
rect 345374 -464 345430 -408
rect 345498 -464 345554 -408
rect 345622 -464 345678 -408
rect 345250 -588 345306 -532
rect 345374 -588 345430 -532
rect 345498 -588 345554 -532
rect 345622 -588 345678 -532
rect 348970 28294 349026 28350
rect 349094 28294 349150 28350
rect 349218 28294 349274 28350
rect 349342 28294 349398 28350
rect 348970 28170 349026 28226
rect 349094 28170 349150 28226
rect 349218 28170 349274 28226
rect 349342 28170 349398 28226
rect 348970 28046 349026 28102
rect 349094 28046 349150 28102
rect 349218 28046 349274 28102
rect 349342 28046 349398 28102
rect 348970 27922 349026 27978
rect 349094 27922 349150 27978
rect 349218 27922 349274 27978
rect 349342 27922 349398 27978
rect 348970 10294 349026 10350
rect 349094 10294 349150 10350
rect 349218 10294 349274 10350
rect 349342 10294 349398 10350
rect 348970 10170 349026 10226
rect 349094 10170 349150 10226
rect 349218 10170 349274 10226
rect 349342 10170 349398 10226
rect 348970 10046 349026 10102
rect 349094 10046 349150 10102
rect 349218 10046 349274 10102
rect 349342 10046 349398 10102
rect 348970 9922 349026 9978
rect 349094 9922 349150 9978
rect 349218 9922 349274 9978
rect 349342 9922 349398 9978
rect 348970 -1176 349026 -1120
rect 349094 -1176 349150 -1120
rect 349218 -1176 349274 -1120
rect 349342 -1176 349398 -1120
rect 348970 -1300 349026 -1244
rect 349094 -1300 349150 -1244
rect 349218 -1300 349274 -1244
rect 349342 -1300 349398 -1244
rect 348970 -1424 349026 -1368
rect 349094 -1424 349150 -1368
rect 349218 -1424 349274 -1368
rect 349342 -1424 349398 -1368
rect 348970 -1548 349026 -1492
rect 349094 -1548 349150 -1492
rect 349218 -1548 349274 -1492
rect 349342 -1548 349398 -1492
rect 363250 22294 363306 22350
rect 363374 22294 363430 22350
rect 363498 22294 363554 22350
rect 363622 22294 363678 22350
rect 363250 22170 363306 22226
rect 363374 22170 363430 22226
rect 363498 22170 363554 22226
rect 363622 22170 363678 22226
rect 363250 22046 363306 22102
rect 363374 22046 363430 22102
rect 363498 22046 363554 22102
rect 363622 22046 363678 22102
rect 363250 21922 363306 21978
rect 363374 21922 363430 21978
rect 363498 21922 363554 21978
rect 363622 21922 363678 21978
rect 363250 4294 363306 4350
rect 363374 4294 363430 4350
rect 363498 4294 363554 4350
rect 363622 4294 363678 4350
rect 363250 4170 363306 4226
rect 363374 4170 363430 4226
rect 363498 4170 363554 4226
rect 363622 4170 363678 4226
rect 363250 4046 363306 4102
rect 363374 4046 363430 4102
rect 363498 4046 363554 4102
rect 363622 4046 363678 4102
rect 363250 3922 363306 3978
rect 363374 3922 363430 3978
rect 363498 3922 363554 3978
rect 363622 3922 363678 3978
rect 363250 -216 363306 -160
rect 363374 -216 363430 -160
rect 363498 -216 363554 -160
rect 363622 -216 363678 -160
rect 363250 -340 363306 -284
rect 363374 -340 363430 -284
rect 363498 -340 363554 -284
rect 363622 -340 363678 -284
rect 363250 -464 363306 -408
rect 363374 -464 363430 -408
rect 363498 -464 363554 -408
rect 363622 -464 363678 -408
rect 363250 -588 363306 -532
rect 363374 -588 363430 -532
rect 363498 -588 363554 -532
rect 363622 -588 363678 -532
rect 366970 28294 367026 28350
rect 367094 28294 367150 28350
rect 367218 28294 367274 28350
rect 367342 28294 367398 28350
rect 366970 28170 367026 28226
rect 367094 28170 367150 28226
rect 367218 28170 367274 28226
rect 367342 28170 367398 28226
rect 366970 28046 367026 28102
rect 367094 28046 367150 28102
rect 367218 28046 367274 28102
rect 367342 28046 367398 28102
rect 366970 27922 367026 27978
rect 367094 27922 367150 27978
rect 367218 27922 367274 27978
rect 367342 27922 367398 27978
rect 366970 10294 367026 10350
rect 367094 10294 367150 10350
rect 367218 10294 367274 10350
rect 367342 10294 367398 10350
rect 366970 10170 367026 10226
rect 367094 10170 367150 10226
rect 367218 10170 367274 10226
rect 367342 10170 367398 10226
rect 366970 10046 367026 10102
rect 367094 10046 367150 10102
rect 367218 10046 367274 10102
rect 367342 10046 367398 10102
rect 366970 9922 367026 9978
rect 367094 9922 367150 9978
rect 367218 9922 367274 9978
rect 367342 9922 367398 9978
rect 366970 -1176 367026 -1120
rect 367094 -1176 367150 -1120
rect 367218 -1176 367274 -1120
rect 367342 -1176 367398 -1120
rect 366970 -1300 367026 -1244
rect 367094 -1300 367150 -1244
rect 367218 -1300 367274 -1244
rect 367342 -1300 367398 -1244
rect 366970 -1424 367026 -1368
rect 367094 -1424 367150 -1368
rect 367218 -1424 367274 -1368
rect 367342 -1424 367398 -1368
rect 366970 -1548 367026 -1492
rect 367094 -1548 367150 -1492
rect 367218 -1548 367274 -1492
rect 367342 -1548 367398 -1492
rect 381250 22294 381306 22350
rect 381374 22294 381430 22350
rect 381498 22294 381554 22350
rect 381622 22294 381678 22350
rect 381250 22170 381306 22226
rect 381374 22170 381430 22226
rect 381498 22170 381554 22226
rect 381622 22170 381678 22226
rect 381250 22046 381306 22102
rect 381374 22046 381430 22102
rect 381498 22046 381554 22102
rect 381622 22046 381678 22102
rect 381250 21922 381306 21978
rect 381374 21922 381430 21978
rect 381498 21922 381554 21978
rect 381622 21922 381678 21978
rect 381250 4294 381306 4350
rect 381374 4294 381430 4350
rect 381498 4294 381554 4350
rect 381622 4294 381678 4350
rect 381250 4170 381306 4226
rect 381374 4170 381430 4226
rect 381498 4170 381554 4226
rect 381622 4170 381678 4226
rect 381250 4046 381306 4102
rect 381374 4046 381430 4102
rect 381498 4046 381554 4102
rect 381622 4046 381678 4102
rect 381250 3922 381306 3978
rect 381374 3922 381430 3978
rect 381498 3922 381554 3978
rect 381622 3922 381678 3978
rect 381250 -216 381306 -160
rect 381374 -216 381430 -160
rect 381498 -216 381554 -160
rect 381622 -216 381678 -160
rect 381250 -340 381306 -284
rect 381374 -340 381430 -284
rect 381498 -340 381554 -284
rect 381622 -340 381678 -284
rect 381250 -464 381306 -408
rect 381374 -464 381430 -408
rect 381498 -464 381554 -408
rect 381622 -464 381678 -408
rect 381250 -588 381306 -532
rect 381374 -588 381430 -532
rect 381498 -588 381554 -532
rect 381622 -588 381678 -532
rect 384970 28294 385026 28350
rect 385094 28294 385150 28350
rect 385218 28294 385274 28350
rect 385342 28294 385398 28350
rect 384970 28170 385026 28226
rect 385094 28170 385150 28226
rect 385218 28170 385274 28226
rect 385342 28170 385398 28226
rect 384970 28046 385026 28102
rect 385094 28046 385150 28102
rect 385218 28046 385274 28102
rect 385342 28046 385398 28102
rect 384970 27922 385026 27978
rect 385094 27922 385150 27978
rect 385218 27922 385274 27978
rect 385342 27922 385398 27978
rect 384970 10294 385026 10350
rect 385094 10294 385150 10350
rect 385218 10294 385274 10350
rect 385342 10294 385398 10350
rect 384970 10170 385026 10226
rect 385094 10170 385150 10226
rect 385218 10170 385274 10226
rect 385342 10170 385398 10226
rect 384970 10046 385026 10102
rect 385094 10046 385150 10102
rect 385218 10046 385274 10102
rect 385342 10046 385398 10102
rect 384970 9922 385026 9978
rect 385094 9922 385150 9978
rect 385218 9922 385274 9978
rect 385342 9922 385398 9978
rect 384970 -1176 385026 -1120
rect 385094 -1176 385150 -1120
rect 385218 -1176 385274 -1120
rect 385342 -1176 385398 -1120
rect 384970 -1300 385026 -1244
rect 385094 -1300 385150 -1244
rect 385218 -1300 385274 -1244
rect 385342 -1300 385398 -1244
rect 384970 -1424 385026 -1368
rect 385094 -1424 385150 -1368
rect 385218 -1424 385274 -1368
rect 385342 -1424 385398 -1368
rect 384970 -1548 385026 -1492
rect 385094 -1548 385150 -1492
rect 385218 -1548 385274 -1492
rect 385342 -1548 385398 -1492
rect 399250 22294 399306 22350
rect 399374 22294 399430 22350
rect 399498 22294 399554 22350
rect 399622 22294 399678 22350
rect 399250 22170 399306 22226
rect 399374 22170 399430 22226
rect 399498 22170 399554 22226
rect 399622 22170 399678 22226
rect 399250 22046 399306 22102
rect 399374 22046 399430 22102
rect 399498 22046 399554 22102
rect 399622 22046 399678 22102
rect 399250 21922 399306 21978
rect 399374 21922 399430 21978
rect 399498 21922 399554 21978
rect 399622 21922 399678 21978
rect 399250 4294 399306 4350
rect 399374 4294 399430 4350
rect 399498 4294 399554 4350
rect 399622 4294 399678 4350
rect 399250 4170 399306 4226
rect 399374 4170 399430 4226
rect 399498 4170 399554 4226
rect 399622 4170 399678 4226
rect 399250 4046 399306 4102
rect 399374 4046 399430 4102
rect 399498 4046 399554 4102
rect 399622 4046 399678 4102
rect 399250 3922 399306 3978
rect 399374 3922 399430 3978
rect 399498 3922 399554 3978
rect 399622 3922 399678 3978
rect 399250 -216 399306 -160
rect 399374 -216 399430 -160
rect 399498 -216 399554 -160
rect 399622 -216 399678 -160
rect 399250 -340 399306 -284
rect 399374 -340 399430 -284
rect 399498 -340 399554 -284
rect 399622 -340 399678 -284
rect 399250 -464 399306 -408
rect 399374 -464 399430 -408
rect 399498 -464 399554 -408
rect 399622 -464 399678 -408
rect 399250 -588 399306 -532
rect 399374 -588 399430 -532
rect 399498 -588 399554 -532
rect 399622 -588 399678 -532
rect 402970 28294 403026 28350
rect 403094 28294 403150 28350
rect 403218 28294 403274 28350
rect 403342 28294 403398 28350
rect 402970 28170 403026 28226
rect 403094 28170 403150 28226
rect 403218 28170 403274 28226
rect 403342 28170 403398 28226
rect 402970 28046 403026 28102
rect 403094 28046 403150 28102
rect 403218 28046 403274 28102
rect 403342 28046 403398 28102
rect 402970 27922 403026 27978
rect 403094 27922 403150 27978
rect 403218 27922 403274 27978
rect 403342 27922 403398 27978
rect 402970 10294 403026 10350
rect 403094 10294 403150 10350
rect 403218 10294 403274 10350
rect 403342 10294 403398 10350
rect 402970 10170 403026 10226
rect 403094 10170 403150 10226
rect 403218 10170 403274 10226
rect 403342 10170 403398 10226
rect 402970 10046 403026 10102
rect 403094 10046 403150 10102
rect 403218 10046 403274 10102
rect 403342 10046 403398 10102
rect 402970 9922 403026 9978
rect 403094 9922 403150 9978
rect 403218 9922 403274 9978
rect 403342 9922 403398 9978
rect 402970 -1176 403026 -1120
rect 403094 -1176 403150 -1120
rect 403218 -1176 403274 -1120
rect 403342 -1176 403398 -1120
rect 402970 -1300 403026 -1244
rect 403094 -1300 403150 -1244
rect 403218 -1300 403274 -1244
rect 403342 -1300 403398 -1244
rect 402970 -1424 403026 -1368
rect 403094 -1424 403150 -1368
rect 403218 -1424 403274 -1368
rect 403342 -1424 403398 -1368
rect 402970 -1548 403026 -1492
rect 403094 -1548 403150 -1492
rect 403218 -1548 403274 -1492
rect 403342 -1548 403398 -1492
rect 417250 22294 417306 22350
rect 417374 22294 417430 22350
rect 417498 22294 417554 22350
rect 417622 22294 417678 22350
rect 417250 22170 417306 22226
rect 417374 22170 417430 22226
rect 417498 22170 417554 22226
rect 417622 22170 417678 22226
rect 417250 22046 417306 22102
rect 417374 22046 417430 22102
rect 417498 22046 417554 22102
rect 417622 22046 417678 22102
rect 417250 21922 417306 21978
rect 417374 21922 417430 21978
rect 417498 21922 417554 21978
rect 417622 21922 417678 21978
rect 417250 4294 417306 4350
rect 417374 4294 417430 4350
rect 417498 4294 417554 4350
rect 417622 4294 417678 4350
rect 417250 4170 417306 4226
rect 417374 4170 417430 4226
rect 417498 4170 417554 4226
rect 417622 4170 417678 4226
rect 417250 4046 417306 4102
rect 417374 4046 417430 4102
rect 417498 4046 417554 4102
rect 417622 4046 417678 4102
rect 417250 3922 417306 3978
rect 417374 3922 417430 3978
rect 417498 3922 417554 3978
rect 417622 3922 417678 3978
rect 417250 -216 417306 -160
rect 417374 -216 417430 -160
rect 417498 -216 417554 -160
rect 417622 -216 417678 -160
rect 417250 -340 417306 -284
rect 417374 -340 417430 -284
rect 417498 -340 417554 -284
rect 417622 -340 417678 -284
rect 417250 -464 417306 -408
rect 417374 -464 417430 -408
rect 417498 -464 417554 -408
rect 417622 -464 417678 -408
rect 417250 -588 417306 -532
rect 417374 -588 417430 -532
rect 417498 -588 417554 -532
rect 417622 -588 417678 -532
rect 420970 28294 421026 28350
rect 421094 28294 421150 28350
rect 421218 28294 421274 28350
rect 421342 28294 421398 28350
rect 420970 28170 421026 28226
rect 421094 28170 421150 28226
rect 421218 28170 421274 28226
rect 421342 28170 421398 28226
rect 420970 28046 421026 28102
rect 421094 28046 421150 28102
rect 421218 28046 421274 28102
rect 421342 28046 421398 28102
rect 420970 27922 421026 27978
rect 421094 27922 421150 27978
rect 421218 27922 421274 27978
rect 421342 27922 421398 27978
rect 420970 10294 421026 10350
rect 421094 10294 421150 10350
rect 421218 10294 421274 10350
rect 421342 10294 421398 10350
rect 420970 10170 421026 10226
rect 421094 10170 421150 10226
rect 421218 10170 421274 10226
rect 421342 10170 421398 10226
rect 420970 10046 421026 10102
rect 421094 10046 421150 10102
rect 421218 10046 421274 10102
rect 421342 10046 421398 10102
rect 420970 9922 421026 9978
rect 421094 9922 421150 9978
rect 421218 9922 421274 9978
rect 421342 9922 421398 9978
rect 420970 -1176 421026 -1120
rect 421094 -1176 421150 -1120
rect 421218 -1176 421274 -1120
rect 421342 -1176 421398 -1120
rect 420970 -1300 421026 -1244
rect 421094 -1300 421150 -1244
rect 421218 -1300 421274 -1244
rect 421342 -1300 421398 -1244
rect 420970 -1424 421026 -1368
rect 421094 -1424 421150 -1368
rect 421218 -1424 421274 -1368
rect 421342 -1424 421398 -1368
rect 420970 -1548 421026 -1492
rect 421094 -1548 421150 -1492
rect 421218 -1548 421274 -1492
rect 421342 -1548 421398 -1492
rect 435250 22294 435306 22350
rect 435374 22294 435430 22350
rect 435498 22294 435554 22350
rect 435622 22294 435678 22350
rect 435250 22170 435306 22226
rect 435374 22170 435430 22226
rect 435498 22170 435554 22226
rect 435622 22170 435678 22226
rect 435250 22046 435306 22102
rect 435374 22046 435430 22102
rect 435498 22046 435554 22102
rect 435622 22046 435678 22102
rect 435250 21922 435306 21978
rect 435374 21922 435430 21978
rect 435498 21922 435554 21978
rect 435622 21922 435678 21978
rect 435250 4294 435306 4350
rect 435374 4294 435430 4350
rect 435498 4294 435554 4350
rect 435622 4294 435678 4350
rect 435250 4170 435306 4226
rect 435374 4170 435430 4226
rect 435498 4170 435554 4226
rect 435622 4170 435678 4226
rect 435250 4046 435306 4102
rect 435374 4046 435430 4102
rect 435498 4046 435554 4102
rect 435622 4046 435678 4102
rect 435250 3922 435306 3978
rect 435374 3922 435430 3978
rect 435498 3922 435554 3978
rect 435622 3922 435678 3978
rect 435250 -216 435306 -160
rect 435374 -216 435430 -160
rect 435498 -216 435554 -160
rect 435622 -216 435678 -160
rect 435250 -340 435306 -284
rect 435374 -340 435430 -284
rect 435498 -340 435554 -284
rect 435622 -340 435678 -284
rect 435250 -464 435306 -408
rect 435374 -464 435430 -408
rect 435498 -464 435554 -408
rect 435622 -464 435678 -408
rect 435250 -588 435306 -532
rect 435374 -588 435430 -532
rect 435498 -588 435554 -532
rect 435622 -588 435678 -532
rect 438970 28294 439026 28350
rect 439094 28294 439150 28350
rect 439218 28294 439274 28350
rect 439342 28294 439398 28350
rect 438970 28170 439026 28226
rect 439094 28170 439150 28226
rect 439218 28170 439274 28226
rect 439342 28170 439398 28226
rect 438970 28046 439026 28102
rect 439094 28046 439150 28102
rect 439218 28046 439274 28102
rect 439342 28046 439398 28102
rect 438970 27922 439026 27978
rect 439094 27922 439150 27978
rect 439218 27922 439274 27978
rect 439342 27922 439398 27978
rect 438970 10294 439026 10350
rect 439094 10294 439150 10350
rect 439218 10294 439274 10350
rect 439342 10294 439398 10350
rect 438970 10170 439026 10226
rect 439094 10170 439150 10226
rect 439218 10170 439274 10226
rect 439342 10170 439398 10226
rect 438970 10046 439026 10102
rect 439094 10046 439150 10102
rect 439218 10046 439274 10102
rect 439342 10046 439398 10102
rect 438970 9922 439026 9978
rect 439094 9922 439150 9978
rect 439218 9922 439274 9978
rect 439342 9922 439398 9978
rect 438970 -1176 439026 -1120
rect 439094 -1176 439150 -1120
rect 439218 -1176 439274 -1120
rect 439342 -1176 439398 -1120
rect 438970 -1300 439026 -1244
rect 439094 -1300 439150 -1244
rect 439218 -1300 439274 -1244
rect 439342 -1300 439398 -1244
rect 438970 -1424 439026 -1368
rect 439094 -1424 439150 -1368
rect 439218 -1424 439274 -1368
rect 439342 -1424 439398 -1368
rect 438970 -1548 439026 -1492
rect 439094 -1548 439150 -1492
rect 439218 -1548 439274 -1492
rect 439342 -1548 439398 -1492
rect 453250 22294 453306 22350
rect 453374 22294 453430 22350
rect 453498 22294 453554 22350
rect 453622 22294 453678 22350
rect 453250 22170 453306 22226
rect 453374 22170 453430 22226
rect 453498 22170 453554 22226
rect 453622 22170 453678 22226
rect 453250 22046 453306 22102
rect 453374 22046 453430 22102
rect 453498 22046 453554 22102
rect 453622 22046 453678 22102
rect 453250 21922 453306 21978
rect 453374 21922 453430 21978
rect 453498 21922 453554 21978
rect 453622 21922 453678 21978
rect 453250 4294 453306 4350
rect 453374 4294 453430 4350
rect 453498 4294 453554 4350
rect 453622 4294 453678 4350
rect 453250 4170 453306 4226
rect 453374 4170 453430 4226
rect 453498 4170 453554 4226
rect 453622 4170 453678 4226
rect 453250 4046 453306 4102
rect 453374 4046 453430 4102
rect 453498 4046 453554 4102
rect 453622 4046 453678 4102
rect 453250 3922 453306 3978
rect 453374 3922 453430 3978
rect 453498 3922 453554 3978
rect 453622 3922 453678 3978
rect 453250 -216 453306 -160
rect 453374 -216 453430 -160
rect 453498 -216 453554 -160
rect 453622 -216 453678 -160
rect 453250 -340 453306 -284
rect 453374 -340 453430 -284
rect 453498 -340 453554 -284
rect 453622 -340 453678 -284
rect 453250 -464 453306 -408
rect 453374 -464 453430 -408
rect 453498 -464 453554 -408
rect 453622 -464 453678 -408
rect 453250 -588 453306 -532
rect 453374 -588 453430 -532
rect 453498 -588 453554 -532
rect 453622 -588 453678 -532
rect 456970 28294 457026 28350
rect 457094 28294 457150 28350
rect 457218 28294 457274 28350
rect 457342 28294 457398 28350
rect 456970 28170 457026 28226
rect 457094 28170 457150 28226
rect 457218 28170 457274 28226
rect 457342 28170 457398 28226
rect 456970 28046 457026 28102
rect 457094 28046 457150 28102
rect 457218 28046 457274 28102
rect 457342 28046 457398 28102
rect 456970 27922 457026 27978
rect 457094 27922 457150 27978
rect 457218 27922 457274 27978
rect 457342 27922 457398 27978
rect 456970 10294 457026 10350
rect 457094 10294 457150 10350
rect 457218 10294 457274 10350
rect 457342 10294 457398 10350
rect 456970 10170 457026 10226
rect 457094 10170 457150 10226
rect 457218 10170 457274 10226
rect 457342 10170 457398 10226
rect 456970 10046 457026 10102
rect 457094 10046 457150 10102
rect 457218 10046 457274 10102
rect 457342 10046 457398 10102
rect 456970 9922 457026 9978
rect 457094 9922 457150 9978
rect 457218 9922 457274 9978
rect 457342 9922 457398 9978
rect 456970 -1176 457026 -1120
rect 457094 -1176 457150 -1120
rect 457218 -1176 457274 -1120
rect 457342 -1176 457398 -1120
rect 456970 -1300 457026 -1244
rect 457094 -1300 457150 -1244
rect 457218 -1300 457274 -1244
rect 457342 -1300 457398 -1244
rect 456970 -1424 457026 -1368
rect 457094 -1424 457150 -1368
rect 457218 -1424 457274 -1368
rect 457342 -1424 457398 -1368
rect 456970 -1548 457026 -1492
rect 457094 -1548 457150 -1492
rect 457218 -1548 457274 -1492
rect 457342 -1548 457398 -1492
rect 471250 22294 471306 22350
rect 471374 22294 471430 22350
rect 471498 22294 471554 22350
rect 471622 22294 471678 22350
rect 471250 22170 471306 22226
rect 471374 22170 471430 22226
rect 471498 22170 471554 22226
rect 471622 22170 471678 22226
rect 471250 22046 471306 22102
rect 471374 22046 471430 22102
rect 471498 22046 471554 22102
rect 471622 22046 471678 22102
rect 471250 21922 471306 21978
rect 471374 21922 471430 21978
rect 471498 21922 471554 21978
rect 471622 21922 471678 21978
rect 471250 4294 471306 4350
rect 471374 4294 471430 4350
rect 471498 4294 471554 4350
rect 471622 4294 471678 4350
rect 471250 4170 471306 4226
rect 471374 4170 471430 4226
rect 471498 4170 471554 4226
rect 471622 4170 471678 4226
rect 471250 4046 471306 4102
rect 471374 4046 471430 4102
rect 471498 4046 471554 4102
rect 471622 4046 471678 4102
rect 471250 3922 471306 3978
rect 471374 3922 471430 3978
rect 471498 3922 471554 3978
rect 471622 3922 471678 3978
rect 471250 -216 471306 -160
rect 471374 -216 471430 -160
rect 471498 -216 471554 -160
rect 471622 -216 471678 -160
rect 471250 -340 471306 -284
rect 471374 -340 471430 -284
rect 471498 -340 471554 -284
rect 471622 -340 471678 -284
rect 471250 -464 471306 -408
rect 471374 -464 471430 -408
rect 471498 -464 471554 -408
rect 471622 -464 471678 -408
rect 471250 -588 471306 -532
rect 471374 -588 471430 -532
rect 471498 -588 471554 -532
rect 471622 -588 471678 -532
rect 474970 28294 475026 28350
rect 475094 28294 475150 28350
rect 475218 28294 475274 28350
rect 475342 28294 475398 28350
rect 474970 28170 475026 28226
rect 475094 28170 475150 28226
rect 475218 28170 475274 28226
rect 475342 28170 475398 28226
rect 474970 28046 475026 28102
rect 475094 28046 475150 28102
rect 475218 28046 475274 28102
rect 475342 28046 475398 28102
rect 474970 27922 475026 27978
rect 475094 27922 475150 27978
rect 475218 27922 475274 27978
rect 475342 27922 475398 27978
rect 474970 10294 475026 10350
rect 475094 10294 475150 10350
rect 475218 10294 475274 10350
rect 475342 10294 475398 10350
rect 474970 10170 475026 10226
rect 475094 10170 475150 10226
rect 475218 10170 475274 10226
rect 475342 10170 475398 10226
rect 474970 10046 475026 10102
rect 475094 10046 475150 10102
rect 475218 10046 475274 10102
rect 475342 10046 475398 10102
rect 474970 9922 475026 9978
rect 475094 9922 475150 9978
rect 475218 9922 475274 9978
rect 475342 9922 475398 9978
rect 474970 -1176 475026 -1120
rect 475094 -1176 475150 -1120
rect 475218 -1176 475274 -1120
rect 475342 -1176 475398 -1120
rect 474970 -1300 475026 -1244
rect 475094 -1300 475150 -1244
rect 475218 -1300 475274 -1244
rect 475342 -1300 475398 -1244
rect 474970 -1424 475026 -1368
rect 475094 -1424 475150 -1368
rect 475218 -1424 475274 -1368
rect 475342 -1424 475398 -1368
rect 474970 -1548 475026 -1492
rect 475094 -1548 475150 -1492
rect 475218 -1548 475274 -1492
rect 475342 -1548 475398 -1492
rect 489250 22294 489306 22350
rect 489374 22294 489430 22350
rect 489498 22294 489554 22350
rect 489622 22294 489678 22350
rect 489250 22170 489306 22226
rect 489374 22170 489430 22226
rect 489498 22170 489554 22226
rect 489622 22170 489678 22226
rect 489250 22046 489306 22102
rect 489374 22046 489430 22102
rect 489498 22046 489554 22102
rect 489622 22046 489678 22102
rect 489250 21922 489306 21978
rect 489374 21922 489430 21978
rect 489498 21922 489554 21978
rect 489622 21922 489678 21978
rect 489250 4294 489306 4350
rect 489374 4294 489430 4350
rect 489498 4294 489554 4350
rect 489622 4294 489678 4350
rect 489250 4170 489306 4226
rect 489374 4170 489430 4226
rect 489498 4170 489554 4226
rect 489622 4170 489678 4226
rect 489250 4046 489306 4102
rect 489374 4046 489430 4102
rect 489498 4046 489554 4102
rect 489622 4046 489678 4102
rect 489250 3922 489306 3978
rect 489374 3922 489430 3978
rect 489498 3922 489554 3978
rect 489622 3922 489678 3978
rect 489250 -216 489306 -160
rect 489374 -216 489430 -160
rect 489498 -216 489554 -160
rect 489622 -216 489678 -160
rect 489250 -340 489306 -284
rect 489374 -340 489430 -284
rect 489498 -340 489554 -284
rect 489622 -340 489678 -284
rect 489250 -464 489306 -408
rect 489374 -464 489430 -408
rect 489498 -464 489554 -408
rect 489622 -464 489678 -408
rect 489250 -588 489306 -532
rect 489374 -588 489430 -532
rect 489498 -588 489554 -532
rect 489622 -588 489678 -532
rect 492970 28294 493026 28350
rect 493094 28294 493150 28350
rect 493218 28294 493274 28350
rect 493342 28294 493398 28350
rect 492970 28170 493026 28226
rect 493094 28170 493150 28226
rect 493218 28170 493274 28226
rect 493342 28170 493398 28226
rect 492970 28046 493026 28102
rect 493094 28046 493150 28102
rect 493218 28046 493274 28102
rect 493342 28046 493398 28102
rect 492970 27922 493026 27978
rect 493094 27922 493150 27978
rect 493218 27922 493274 27978
rect 493342 27922 493398 27978
rect 492970 10294 493026 10350
rect 493094 10294 493150 10350
rect 493218 10294 493274 10350
rect 493342 10294 493398 10350
rect 492970 10170 493026 10226
rect 493094 10170 493150 10226
rect 493218 10170 493274 10226
rect 493342 10170 493398 10226
rect 492970 10046 493026 10102
rect 493094 10046 493150 10102
rect 493218 10046 493274 10102
rect 493342 10046 493398 10102
rect 492970 9922 493026 9978
rect 493094 9922 493150 9978
rect 493218 9922 493274 9978
rect 493342 9922 493398 9978
rect 492970 -1176 493026 -1120
rect 493094 -1176 493150 -1120
rect 493218 -1176 493274 -1120
rect 493342 -1176 493398 -1120
rect 492970 -1300 493026 -1244
rect 493094 -1300 493150 -1244
rect 493218 -1300 493274 -1244
rect 493342 -1300 493398 -1244
rect 492970 -1424 493026 -1368
rect 493094 -1424 493150 -1368
rect 493218 -1424 493274 -1368
rect 493342 -1424 493398 -1368
rect 492970 -1548 493026 -1492
rect 493094 -1548 493150 -1492
rect 493218 -1548 493274 -1492
rect 493342 -1548 493398 -1492
rect 507250 22294 507306 22350
rect 507374 22294 507430 22350
rect 507498 22294 507554 22350
rect 507622 22294 507678 22350
rect 507250 22170 507306 22226
rect 507374 22170 507430 22226
rect 507498 22170 507554 22226
rect 507622 22170 507678 22226
rect 507250 22046 507306 22102
rect 507374 22046 507430 22102
rect 507498 22046 507554 22102
rect 507622 22046 507678 22102
rect 507250 21922 507306 21978
rect 507374 21922 507430 21978
rect 507498 21922 507554 21978
rect 507622 21922 507678 21978
rect 507250 4294 507306 4350
rect 507374 4294 507430 4350
rect 507498 4294 507554 4350
rect 507622 4294 507678 4350
rect 507250 4170 507306 4226
rect 507374 4170 507430 4226
rect 507498 4170 507554 4226
rect 507622 4170 507678 4226
rect 507250 4046 507306 4102
rect 507374 4046 507430 4102
rect 507498 4046 507554 4102
rect 507622 4046 507678 4102
rect 507250 3922 507306 3978
rect 507374 3922 507430 3978
rect 507498 3922 507554 3978
rect 507622 3922 507678 3978
rect 507250 -216 507306 -160
rect 507374 -216 507430 -160
rect 507498 -216 507554 -160
rect 507622 -216 507678 -160
rect 507250 -340 507306 -284
rect 507374 -340 507430 -284
rect 507498 -340 507554 -284
rect 507622 -340 507678 -284
rect 507250 -464 507306 -408
rect 507374 -464 507430 -408
rect 507498 -464 507554 -408
rect 507622 -464 507678 -408
rect 507250 -588 507306 -532
rect 507374 -588 507430 -532
rect 507498 -588 507554 -532
rect 507622 -588 507678 -532
rect 510970 28294 511026 28350
rect 511094 28294 511150 28350
rect 511218 28294 511274 28350
rect 511342 28294 511398 28350
rect 510970 28170 511026 28226
rect 511094 28170 511150 28226
rect 511218 28170 511274 28226
rect 511342 28170 511398 28226
rect 510970 28046 511026 28102
rect 511094 28046 511150 28102
rect 511218 28046 511274 28102
rect 511342 28046 511398 28102
rect 510970 27922 511026 27978
rect 511094 27922 511150 27978
rect 511218 27922 511274 27978
rect 511342 27922 511398 27978
rect 510970 10294 511026 10350
rect 511094 10294 511150 10350
rect 511218 10294 511274 10350
rect 511342 10294 511398 10350
rect 510970 10170 511026 10226
rect 511094 10170 511150 10226
rect 511218 10170 511274 10226
rect 511342 10170 511398 10226
rect 510970 10046 511026 10102
rect 511094 10046 511150 10102
rect 511218 10046 511274 10102
rect 511342 10046 511398 10102
rect 510970 9922 511026 9978
rect 511094 9922 511150 9978
rect 511218 9922 511274 9978
rect 511342 9922 511398 9978
rect 510970 -1176 511026 -1120
rect 511094 -1176 511150 -1120
rect 511218 -1176 511274 -1120
rect 511342 -1176 511398 -1120
rect 510970 -1300 511026 -1244
rect 511094 -1300 511150 -1244
rect 511218 -1300 511274 -1244
rect 511342 -1300 511398 -1244
rect 510970 -1424 511026 -1368
rect 511094 -1424 511150 -1368
rect 511218 -1424 511274 -1368
rect 511342 -1424 511398 -1368
rect 510970 -1548 511026 -1492
rect 511094 -1548 511150 -1492
rect 511218 -1548 511274 -1492
rect 511342 -1548 511398 -1492
rect 525250 22294 525306 22350
rect 525374 22294 525430 22350
rect 525498 22294 525554 22350
rect 525622 22294 525678 22350
rect 525250 22170 525306 22226
rect 525374 22170 525430 22226
rect 525498 22170 525554 22226
rect 525622 22170 525678 22226
rect 525250 22046 525306 22102
rect 525374 22046 525430 22102
rect 525498 22046 525554 22102
rect 525622 22046 525678 22102
rect 525250 21922 525306 21978
rect 525374 21922 525430 21978
rect 525498 21922 525554 21978
rect 525622 21922 525678 21978
rect 525250 4294 525306 4350
rect 525374 4294 525430 4350
rect 525498 4294 525554 4350
rect 525622 4294 525678 4350
rect 525250 4170 525306 4226
rect 525374 4170 525430 4226
rect 525498 4170 525554 4226
rect 525622 4170 525678 4226
rect 525250 4046 525306 4102
rect 525374 4046 525430 4102
rect 525498 4046 525554 4102
rect 525622 4046 525678 4102
rect 525250 3922 525306 3978
rect 525374 3922 525430 3978
rect 525498 3922 525554 3978
rect 525622 3922 525678 3978
rect 525250 -216 525306 -160
rect 525374 -216 525430 -160
rect 525498 -216 525554 -160
rect 525622 -216 525678 -160
rect 525250 -340 525306 -284
rect 525374 -340 525430 -284
rect 525498 -340 525554 -284
rect 525622 -340 525678 -284
rect 525250 -464 525306 -408
rect 525374 -464 525430 -408
rect 525498 -464 525554 -408
rect 525622 -464 525678 -408
rect 525250 -588 525306 -532
rect 525374 -588 525430 -532
rect 525498 -588 525554 -532
rect 525622 -588 525678 -532
rect 528970 28294 529026 28350
rect 529094 28294 529150 28350
rect 529218 28294 529274 28350
rect 529342 28294 529398 28350
rect 528970 28170 529026 28226
rect 529094 28170 529150 28226
rect 529218 28170 529274 28226
rect 529342 28170 529398 28226
rect 528970 28046 529026 28102
rect 529094 28046 529150 28102
rect 529218 28046 529274 28102
rect 529342 28046 529398 28102
rect 528970 27922 529026 27978
rect 529094 27922 529150 27978
rect 529218 27922 529274 27978
rect 529342 27922 529398 27978
rect 528970 10294 529026 10350
rect 529094 10294 529150 10350
rect 529218 10294 529274 10350
rect 529342 10294 529398 10350
rect 528970 10170 529026 10226
rect 529094 10170 529150 10226
rect 529218 10170 529274 10226
rect 529342 10170 529398 10226
rect 528970 10046 529026 10102
rect 529094 10046 529150 10102
rect 529218 10046 529274 10102
rect 529342 10046 529398 10102
rect 528970 9922 529026 9978
rect 529094 9922 529150 9978
rect 529218 9922 529274 9978
rect 529342 9922 529398 9978
rect 528970 -1176 529026 -1120
rect 529094 -1176 529150 -1120
rect 529218 -1176 529274 -1120
rect 529342 -1176 529398 -1120
rect 528970 -1300 529026 -1244
rect 529094 -1300 529150 -1244
rect 529218 -1300 529274 -1244
rect 529342 -1300 529398 -1244
rect 528970 -1424 529026 -1368
rect 529094 -1424 529150 -1368
rect 529218 -1424 529274 -1368
rect 529342 -1424 529398 -1368
rect 528970 -1548 529026 -1492
rect 529094 -1548 529150 -1492
rect 529218 -1548 529274 -1492
rect 529342 -1548 529398 -1492
rect 543250 22294 543306 22350
rect 543374 22294 543430 22350
rect 543498 22294 543554 22350
rect 543622 22294 543678 22350
rect 543250 22170 543306 22226
rect 543374 22170 543430 22226
rect 543498 22170 543554 22226
rect 543622 22170 543678 22226
rect 543250 22046 543306 22102
rect 543374 22046 543430 22102
rect 543498 22046 543554 22102
rect 543622 22046 543678 22102
rect 543250 21922 543306 21978
rect 543374 21922 543430 21978
rect 543498 21922 543554 21978
rect 543622 21922 543678 21978
rect 543250 4294 543306 4350
rect 543374 4294 543430 4350
rect 543498 4294 543554 4350
rect 543622 4294 543678 4350
rect 543250 4170 543306 4226
rect 543374 4170 543430 4226
rect 543498 4170 543554 4226
rect 543622 4170 543678 4226
rect 543250 4046 543306 4102
rect 543374 4046 543430 4102
rect 543498 4046 543554 4102
rect 543622 4046 543678 4102
rect 543250 3922 543306 3978
rect 543374 3922 543430 3978
rect 543498 3922 543554 3978
rect 543622 3922 543678 3978
rect 543250 -216 543306 -160
rect 543374 -216 543430 -160
rect 543498 -216 543554 -160
rect 543622 -216 543678 -160
rect 543250 -340 543306 -284
rect 543374 -340 543430 -284
rect 543498 -340 543554 -284
rect 543622 -340 543678 -284
rect 543250 -464 543306 -408
rect 543374 -464 543430 -408
rect 543498 -464 543554 -408
rect 543622 -464 543678 -408
rect 543250 -588 543306 -532
rect 543374 -588 543430 -532
rect 543498 -588 543554 -532
rect 543622 -588 543678 -532
rect 546970 28294 547026 28350
rect 547094 28294 547150 28350
rect 547218 28294 547274 28350
rect 547342 28294 547398 28350
rect 546970 28170 547026 28226
rect 547094 28170 547150 28226
rect 547218 28170 547274 28226
rect 547342 28170 547398 28226
rect 546970 28046 547026 28102
rect 547094 28046 547150 28102
rect 547218 28046 547274 28102
rect 547342 28046 547398 28102
rect 546970 27922 547026 27978
rect 547094 27922 547150 27978
rect 547218 27922 547274 27978
rect 547342 27922 547398 27978
rect 546970 10294 547026 10350
rect 547094 10294 547150 10350
rect 547218 10294 547274 10350
rect 547342 10294 547398 10350
rect 546970 10170 547026 10226
rect 547094 10170 547150 10226
rect 547218 10170 547274 10226
rect 547342 10170 547398 10226
rect 546970 10046 547026 10102
rect 547094 10046 547150 10102
rect 547218 10046 547274 10102
rect 547342 10046 547398 10102
rect 546970 9922 547026 9978
rect 547094 9922 547150 9978
rect 547218 9922 547274 9978
rect 547342 9922 547398 9978
rect 546970 -1176 547026 -1120
rect 547094 -1176 547150 -1120
rect 547218 -1176 547274 -1120
rect 547342 -1176 547398 -1120
rect 546970 -1300 547026 -1244
rect 547094 -1300 547150 -1244
rect 547218 -1300 547274 -1244
rect 547342 -1300 547398 -1244
rect 546970 -1424 547026 -1368
rect 547094 -1424 547150 -1368
rect 547218 -1424 547274 -1368
rect 547342 -1424 547398 -1368
rect 546970 -1548 547026 -1492
rect 547094 -1548 547150 -1492
rect 547218 -1548 547274 -1492
rect 547342 -1548 547398 -1492
rect 561250 22294 561306 22350
rect 561374 22294 561430 22350
rect 561498 22294 561554 22350
rect 561622 22294 561678 22350
rect 561250 22170 561306 22226
rect 561374 22170 561430 22226
rect 561498 22170 561554 22226
rect 561622 22170 561678 22226
rect 561250 22046 561306 22102
rect 561374 22046 561430 22102
rect 561498 22046 561554 22102
rect 561622 22046 561678 22102
rect 561250 21922 561306 21978
rect 561374 21922 561430 21978
rect 561498 21922 561554 21978
rect 561622 21922 561678 21978
rect 561250 4294 561306 4350
rect 561374 4294 561430 4350
rect 561498 4294 561554 4350
rect 561622 4294 561678 4350
rect 561250 4170 561306 4226
rect 561374 4170 561430 4226
rect 561498 4170 561554 4226
rect 561622 4170 561678 4226
rect 561250 4046 561306 4102
rect 561374 4046 561430 4102
rect 561498 4046 561554 4102
rect 561622 4046 561678 4102
rect 561250 3922 561306 3978
rect 561374 3922 561430 3978
rect 561498 3922 561554 3978
rect 561622 3922 561678 3978
rect 561250 -216 561306 -160
rect 561374 -216 561430 -160
rect 561498 -216 561554 -160
rect 561622 -216 561678 -160
rect 561250 -340 561306 -284
rect 561374 -340 561430 -284
rect 561498 -340 561554 -284
rect 561622 -340 561678 -284
rect 561250 -464 561306 -408
rect 561374 -464 561430 -408
rect 561498 -464 561554 -408
rect 561622 -464 561678 -408
rect 561250 -588 561306 -532
rect 561374 -588 561430 -532
rect 561498 -588 561554 -532
rect 561622 -588 561678 -532
rect 564970 598116 565026 598172
rect 565094 598116 565150 598172
rect 565218 598116 565274 598172
rect 565342 598116 565398 598172
rect 564970 597992 565026 598048
rect 565094 597992 565150 598048
rect 565218 597992 565274 598048
rect 565342 597992 565398 598048
rect 564970 597868 565026 597924
rect 565094 597868 565150 597924
rect 565218 597868 565274 597924
rect 565342 597868 565398 597924
rect 564970 597744 565026 597800
rect 565094 597744 565150 597800
rect 565218 597744 565274 597800
rect 565342 597744 565398 597800
rect 564970 586294 565026 586350
rect 565094 586294 565150 586350
rect 565218 586294 565274 586350
rect 565342 586294 565398 586350
rect 564970 586170 565026 586226
rect 565094 586170 565150 586226
rect 565218 586170 565274 586226
rect 565342 586170 565398 586226
rect 564970 586046 565026 586102
rect 565094 586046 565150 586102
rect 565218 586046 565274 586102
rect 565342 586046 565398 586102
rect 564970 585922 565026 585978
rect 565094 585922 565150 585978
rect 565218 585922 565274 585978
rect 565342 585922 565398 585978
rect 564970 568294 565026 568350
rect 565094 568294 565150 568350
rect 565218 568294 565274 568350
rect 565342 568294 565398 568350
rect 564970 568170 565026 568226
rect 565094 568170 565150 568226
rect 565218 568170 565274 568226
rect 565342 568170 565398 568226
rect 564970 568046 565026 568102
rect 565094 568046 565150 568102
rect 565218 568046 565274 568102
rect 565342 568046 565398 568102
rect 564970 567922 565026 567978
rect 565094 567922 565150 567978
rect 565218 567922 565274 567978
rect 565342 567922 565398 567978
rect 564970 550294 565026 550350
rect 565094 550294 565150 550350
rect 565218 550294 565274 550350
rect 565342 550294 565398 550350
rect 564970 550170 565026 550226
rect 565094 550170 565150 550226
rect 565218 550170 565274 550226
rect 565342 550170 565398 550226
rect 564970 550046 565026 550102
rect 565094 550046 565150 550102
rect 565218 550046 565274 550102
rect 565342 550046 565398 550102
rect 564970 549922 565026 549978
rect 565094 549922 565150 549978
rect 565218 549922 565274 549978
rect 565342 549922 565398 549978
rect 564970 532294 565026 532350
rect 565094 532294 565150 532350
rect 565218 532294 565274 532350
rect 565342 532294 565398 532350
rect 564970 532170 565026 532226
rect 565094 532170 565150 532226
rect 565218 532170 565274 532226
rect 565342 532170 565398 532226
rect 564970 532046 565026 532102
rect 565094 532046 565150 532102
rect 565218 532046 565274 532102
rect 565342 532046 565398 532102
rect 564970 531922 565026 531978
rect 565094 531922 565150 531978
rect 565218 531922 565274 531978
rect 565342 531922 565398 531978
rect 564970 514294 565026 514350
rect 565094 514294 565150 514350
rect 565218 514294 565274 514350
rect 565342 514294 565398 514350
rect 564970 514170 565026 514226
rect 565094 514170 565150 514226
rect 565218 514170 565274 514226
rect 565342 514170 565398 514226
rect 564970 514046 565026 514102
rect 565094 514046 565150 514102
rect 565218 514046 565274 514102
rect 565342 514046 565398 514102
rect 564970 513922 565026 513978
rect 565094 513922 565150 513978
rect 565218 513922 565274 513978
rect 565342 513922 565398 513978
rect 564970 496294 565026 496350
rect 565094 496294 565150 496350
rect 565218 496294 565274 496350
rect 565342 496294 565398 496350
rect 564970 496170 565026 496226
rect 565094 496170 565150 496226
rect 565218 496170 565274 496226
rect 565342 496170 565398 496226
rect 564970 496046 565026 496102
rect 565094 496046 565150 496102
rect 565218 496046 565274 496102
rect 565342 496046 565398 496102
rect 564970 495922 565026 495978
rect 565094 495922 565150 495978
rect 565218 495922 565274 495978
rect 565342 495922 565398 495978
rect 564970 478294 565026 478350
rect 565094 478294 565150 478350
rect 565218 478294 565274 478350
rect 565342 478294 565398 478350
rect 564970 478170 565026 478226
rect 565094 478170 565150 478226
rect 565218 478170 565274 478226
rect 565342 478170 565398 478226
rect 564970 478046 565026 478102
rect 565094 478046 565150 478102
rect 565218 478046 565274 478102
rect 565342 478046 565398 478102
rect 564970 477922 565026 477978
rect 565094 477922 565150 477978
rect 565218 477922 565274 477978
rect 565342 477922 565398 477978
rect 564970 460294 565026 460350
rect 565094 460294 565150 460350
rect 565218 460294 565274 460350
rect 565342 460294 565398 460350
rect 564970 460170 565026 460226
rect 565094 460170 565150 460226
rect 565218 460170 565274 460226
rect 565342 460170 565398 460226
rect 564970 460046 565026 460102
rect 565094 460046 565150 460102
rect 565218 460046 565274 460102
rect 565342 460046 565398 460102
rect 564970 459922 565026 459978
rect 565094 459922 565150 459978
rect 565218 459922 565274 459978
rect 565342 459922 565398 459978
rect 564970 442294 565026 442350
rect 565094 442294 565150 442350
rect 565218 442294 565274 442350
rect 565342 442294 565398 442350
rect 564970 442170 565026 442226
rect 565094 442170 565150 442226
rect 565218 442170 565274 442226
rect 565342 442170 565398 442226
rect 564970 442046 565026 442102
rect 565094 442046 565150 442102
rect 565218 442046 565274 442102
rect 565342 442046 565398 442102
rect 564970 441922 565026 441978
rect 565094 441922 565150 441978
rect 565218 441922 565274 441978
rect 565342 441922 565398 441978
rect 564970 424294 565026 424350
rect 565094 424294 565150 424350
rect 565218 424294 565274 424350
rect 565342 424294 565398 424350
rect 564970 424170 565026 424226
rect 565094 424170 565150 424226
rect 565218 424170 565274 424226
rect 565342 424170 565398 424226
rect 564970 424046 565026 424102
rect 565094 424046 565150 424102
rect 565218 424046 565274 424102
rect 565342 424046 565398 424102
rect 564970 423922 565026 423978
rect 565094 423922 565150 423978
rect 565218 423922 565274 423978
rect 565342 423922 565398 423978
rect 564970 406294 565026 406350
rect 565094 406294 565150 406350
rect 565218 406294 565274 406350
rect 565342 406294 565398 406350
rect 564970 406170 565026 406226
rect 565094 406170 565150 406226
rect 565218 406170 565274 406226
rect 565342 406170 565398 406226
rect 564970 406046 565026 406102
rect 565094 406046 565150 406102
rect 565218 406046 565274 406102
rect 565342 406046 565398 406102
rect 564970 405922 565026 405978
rect 565094 405922 565150 405978
rect 565218 405922 565274 405978
rect 565342 405922 565398 405978
rect 564970 388294 565026 388350
rect 565094 388294 565150 388350
rect 565218 388294 565274 388350
rect 565342 388294 565398 388350
rect 564970 388170 565026 388226
rect 565094 388170 565150 388226
rect 565218 388170 565274 388226
rect 565342 388170 565398 388226
rect 564970 388046 565026 388102
rect 565094 388046 565150 388102
rect 565218 388046 565274 388102
rect 565342 388046 565398 388102
rect 564970 387922 565026 387978
rect 565094 387922 565150 387978
rect 565218 387922 565274 387978
rect 565342 387922 565398 387978
rect 564970 370294 565026 370350
rect 565094 370294 565150 370350
rect 565218 370294 565274 370350
rect 565342 370294 565398 370350
rect 564970 370170 565026 370226
rect 565094 370170 565150 370226
rect 565218 370170 565274 370226
rect 565342 370170 565398 370226
rect 564970 370046 565026 370102
rect 565094 370046 565150 370102
rect 565218 370046 565274 370102
rect 565342 370046 565398 370102
rect 564970 369922 565026 369978
rect 565094 369922 565150 369978
rect 565218 369922 565274 369978
rect 565342 369922 565398 369978
rect 564970 352294 565026 352350
rect 565094 352294 565150 352350
rect 565218 352294 565274 352350
rect 565342 352294 565398 352350
rect 564970 352170 565026 352226
rect 565094 352170 565150 352226
rect 565218 352170 565274 352226
rect 565342 352170 565398 352226
rect 564970 352046 565026 352102
rect 565094 352046 565150 352102
rect 565218 352046 565274 352102
rect 565342 352046 565398 352102
rect 564970 351922 565026 351978
rect 565094 351922 565150 351978
rect 565218 351922 565274 351978
rect 565342 351922 565398 351978
rect 564970 334294 565026 334350
rect 565094 334294 565150 334350
rect 565218 334294 565274 334350
rect 565342 334294 565398 334350
rect 564970 334170 565026 334226
rect 565094 334170 565150 334226
rect 565218 334170 565274 334226
rect 565342 334170 565398 334226
rect 564970 334046 565026 334102
rect 565094 334046 565150 334102
rect 565218 334046 565274 334102
rect 565342 334046 565398 334102
rect 564970 333922 565026 333978
rect 565094 333922 565150 333978
rect 565218 333922 565274 333978
rect 565342 333922 565398 333978
rect 564970 316294 565026 316350
rect 565094 316294 565150 316350
rect 565218 316294 565274 316350
rect 565342 316294 565398 316350
rect 564970 316170 565026 316226
rect 565094 316170 565150 316226
rect 565218 316170 565274 316226
rect 565342 316170 565398 316226
rect 564970 316046 565026 316102
rect 565094 316046 565150 316102
rect 565218 316046 565274 316102
rect 565342 316046 565398 316102
rect 564970 315922 565026 315978
rect 565094 315922 565150 315978
rect 565218 315922 565274 315978
rect 565342 315922 565398 315978
rect 564970 298294 565026 298350
rect 565094 298294 565150 298350
rect 565218 298294 565274 298350
rect 565342 298294 565398 298350
rect 564970 298170 565026 298226
rect 565094 298170 565150 298226
rect 565218 298170 565274 298226
rect 565342 298170 565398 298226
rect 564970 298046 565026 298102
rect 565094 298046 565150 298102
rect 565218 298046 565274 298102
rect 565342 298046 565398 298102
rect 564970 297922 565026 297978
rect 565094 297922 565150 297978
rect 565218 297922 565274 297978
rect 565342 297922 565398 297978
rect 564970 280294 565026 280350
rect 565094 280294 565150 280350
rect 565218 280294 565274 280350
rect 565342 280294 565398 280350
rect 564970 280170 565026 280226
rect 565094 280170 565150 280226
rect 565218 280170 565274 280226
rect 565342 280170 565398 280226
rect 564970 280046 565026 280102
rect 565094 280046 565150 280102
rect 565218 280046 565274 280102
rect 565342 280046 565398 280102
rect 564970 279922 565026 279978
rect 565094 279922 565150 279978
rect 565218 279922 565274 279978
rect 565342 279922 565398 279978
rect 564970 262294 565026 262350
rect 565094 262294 565150 262350
rect 565218 262294 565274 262350
rect 565342 262294 565398 262350
rect 564970 262170 565026 262226
rect 565094 262170 565150 262226
rect 565218 262170 565274 262226
rect 565342 262170 565398 262226
rect 564970 262046 565026 262102
rect 565094 262046 565150 262102
rect 565218 262046 565274 262102
rect 565342 262046 565398 262102
rect 564970 261922 565026 261978
rect 565094 261922 565150 261978
rect 565218 261922 565274 261978
rect 565342 261922 565398 261978
rect 564970 244294 565026 244350
rect 565094 244294 565150 244350
rect 565218 244294 565274 244350
rect 565342 244294 565398 244350
rect 564970 244170 565026 244226
rect 565094 244170 565150 244226
rect 565218 244170 565274 244226
rect 565342 244170 565398 244226
rect 564970 244046 565026 244102
rect 565094 244046 565150 244102
rect 565218 244046 565274 244102
rect 565342 244046 565398 244102
rect 564970 243922 565026 243978
rect 565094 243922 565150 243978
rect 565218 243922 565274 243978
rect 565342 243922 565398 243978
rect 564970 226294 565026 226350
rect 565094 226294 565150 226350
rect 565218 226294 565274 226350
rect 565342 226294 565398 226350
rect 564970 226170 565026 226226
rect 565094 226170 565150 226226
rect 565218 226170 565274 226226
rect 565342 226170 565398 226226
rect 564970 226046 565026 226102
rect 565094 226046 565150 226102
rect 565218 226046 565274 226102
rect 565342 226046 565398 226102
rect 564970 225922 565026 225978
rect 565094 225922 565150 225978
rect 565218 225922 565274 225978
rect 565342 225922 565398 225978
rect 564970 208294 565026 208350
rect 565094 208294 565150 208350
rect 565218 208294 565274 208350
rect 565342 208294 565398 208350
rect 564970 208170 565026 208226
rect 565094 208170 565150 208226
rect 565218 208170 565274 208226
rect 565342 208170 565398 208226
rect 564970 208046 565026 208102
rect 565094 208046 565150 208102
rect 565218 208046 565274 208102
rect 565342 208046 565398 208102
rect 564970 207922 565026 207978
rect 565094 207922 565150 207978
rect 565218 207922 565274 207978
rect 565342 207922 565398 207978
rect 564970 190294 565026 190350
rect 565094 190294 565150 190350
rect 565218 190294 565274 190350
rect 565342 190294 565398 190350
rect 564970 190170 565026 190226
rect 565094 190170 565150 190226
rect 565218 190170 565274 190226
rect 565342 190170 565398 190226
rect 564970 190046 565026 190102
rect 565094 190046 565150 190102
rect 565218 190046 565274 190102
rect 565342 190046 565398 190102
rect 564970 189922 565026 189978
rect 565094 189922 565150 189978
rect 565218 189922 565274 189978
rect 565342 189922 565398 189978
rect 564970 172294 565026 172350
rect 565094 172294 565150 172350
rect 565218 172294 565274 172350
rect 565342 172294 565398 172350
rect 564970 172170 565026 172226
rect 565094 172170 565150 172226
rect 565218 172170 565274 172226
rect 565342 172170 565398 172226
rect 564970 172046 565026 172102
rect 565094 172046 565150 172102
rect 565218 172046 565274 172102
rect 565342 172046 565398 172102
rect 564970 171922 565026 171978
rect 565094 171922 565150 171978
rect 565218 171922 565274 171978
rect 565342 171922 565398 171978
rect 564970 154294 565026 154350
rect 565094 154294 565150 154350
rect 565218 154294 565274 154350
rect 565342 154294 565398 154350
rect 564970 154170 565026 154226
rect 565094 154170 565150 154226
rect 565218 154170 565274 154226
rect 565342 154170 565398 154226
rect 564970 154046 565026 154102
rect 565094 154046 565150 154102
rect 565218 154046 565274 154102
rect 565342 154046 565398 154102
rect 564970 153922 565026 153978
rect 565094 153922 565150 153978
rect 565218 153922 565274 153978
rect 565342 153922 565398 153978
rect 564970 136294 565026 136350
rect 565094 136294 565150 136350
rect 565218 136294 565274 136350
rect 565342 136294 565398 136350
rect 564970 136170 565026 136226
rect 565094 136170 565150 136226
rect 565218 136170 565274 136226
rect 565342 136170 565398 136226
rect 564970 136046 565026 136102
rect 565094 136046 565150 136102
rect 565218 136046 565274 136102
rect 565342 136046 565398 136102
rect 564970 135922 565026 135978
rect 565094 135922 565150 135978
rect 565218 135922 565274 135978
rect 565342 135922 565398 135978
rect 564970 118294 565026 118350
rect 565094 118294 565150 118350
rect 565218 118294 565274 118350
rect 565342 118294 565398 118350
rect 564970 118170 565026 118226
rect 565094 118170 565150 118226
rect 565218 118170 565274 118226
rect 565342 118170 565398 118226
rect 564970 118046 565026 118102
rect 565094 118046 565150 118102
rect 565218 118046 565274 118102
rect 565342 118046 565398 118102
rect 564970 117922 565026 117978
rect 565094 117922 565150 117978
rect 565218 117922 565274 117978
rect 565342 117922 565398 117978
rect 564970 100294 565026 100350
rect 565094 100294 565150 100350
rect 565218 100294 565274 100350
rect 565342 100294 565398 100350
rect 564970 100170 565026 100226
rect 565094 100170 565150 100226
rect 565218 100170 565274 100226
rect 565342 100170 565398 100226
rect 564970 100046 565026 100102
rect 565094 100046 565150 100102
rect 565218 100046 565274 100102
rect 565342 100046 565398 100102
rect 564970 99922 565026 99978
rect 565094 99922 565150 99978
rect 565218 99922 565274 99978
rect 565342 99922 565398 99978
rect 564970 82294 565026 82350
rect 565094 82294 565150 82350
rect 565218 82294 565274 82350
rect 565342 82294 565398 82350
rect 564970 82170 565026 82226
rect 565094 82170 565150 82226
rect 565218 82170 565274 82226
rect 565342 82170 565398 82226
rect 564970 82046 565026 82102
rect 565094 82046 565150 82102
rect 565218 82046 565274 82102
rect 565342 82046 565398 82102
rect 564970 81922 565026 81978
rect 565094 81922 565150 81978
rect 565218 81922 565274 81978
rect 565342 81922 565398 81978
rect 564970 64294 565026 64350
rect 565094 64294 565150 64350
rect 565218 64294 565274 64350
rect 565342 64294 565398 64350
rect 564970 64170 565026 64226
rect 565094 64170 565150 64226
rect 565218 64170 565274 64226
rect 565342 64170 565398 64226
rect 564970 64046 565026 64102
rect 565094 64046 565150 64102
rect 565218 64046 565274 64102
rect 565342 64046 565398 64102
rect 564970 63922 565026 63978
rect 565094 63922 565150 63978
rect 565218 63922 565274 63978
rect 565342 63922 565398 63978
rect 564970 46294 565026 46350
rect 565094 46294 565150 46350
rect 565218 46294 565274 46350
rect 565342 46294 565398 46350
rect 564970 46170 565026 46226
rect 565094 46170 565150 46226
rect 565218 46170 565274 46226
rect 565342 46170 565398 46226
rect 564970 46046 565026 46102
rect 565094 46046 565150 46102
rect 565218 46046 565274 46102
rect 565342 46046 565398 46102
rect 564970 45922 565026 45978
rect 565094 45922 565150 45978
rect 565218 45922 565274 45978
rect 565342 45922 565398 45978
rect 564970 28294 565026 28350
rect 565094 28294 565150 28350
rect 565218 28294 565274 28350
rect 565342 28294 565398 28350
rect 564970 28170 565026 28226
rect 565094 28170 565150 28226
rect 565218 28170 565274 28226
rect 565342 28170 565398 28226
rect 564970 28046 565026 28102
rect 565094 28046 565150 28102
rect 565218 28046 565274 28102
rect 565342 28046 565398 28102
rect 564970 27922 565026 27978
rect 565094 27922 565150 27978
rect 565218 27922 565274 27978
rect 565342 27922 565398 27978
rect 564970 10294 565026 10350
rect 565094 10294 565150 10350
rect 565218 10294 565274 10350
rect 565342 10294 565398 10350
rect 564970 10170 565026 10226
rect 565094 10170 565150 10226
rect 565218 10170 565274 10226
rect 565342 10170 565398 10226
rect 564970 10046 565026 10102
rect 565094 10046 565150 10102
rect 565218 10046 565274 10102
rect 565342 10046 565398 10102
rect 564970 9922 565026 9978
rect 565094 9922 565150 9978
rect 565218 9922 565274 9978
rect 565342 9922 565398 9978
rect 564970 -1176 565026 -1120
rect 565094 -1176 565150 -1120
rect 565218 -1176 565274 -1120
rect 565342 -1176 565398 -1120
rect 564970 -1300 565026 -1244
rect 565094 -1300 565150 -1244
rect 565218 -1300 565274 -1244
rect 565342 -1300 565398 -1244
rect 564970 -1424 565026 -1368
rect 565094 -1424 565150 -1368
rect 565218 -1424 565274 -1368
rect 565342 -1424 565398 -1368
rect 564970 -1548 565026 -1492
rect 565094 -1548 565150 -1492
rect 565218 -1548 565274 -1492
rect 565342 -1548 565398 -1492
rect 579250 597156 579306 597212
rect 579374 597156 579430 597212
rect 579498 597156 579554 597212
rect 579622 597156 579678 597212
rect 579250 597032 579306 597088
rect 579374 597032 579430 597088
rect 579498 597032 579554 597088
rect 579622 597032 579678 597088
rect 579250 596908 579306 596964
rect 579374 596908 579430 596964
rect 579498 596908 579554 596964
rect 579622 596908 579678 596964
rect 579250 596784 579306 596840
rect 579374 596784 579430 596840
rect 579498 596784 579554 596840
rect 579622 596784 579678 596840
rect 579250 580294 579306 580350
rect 579374 580294 579430 580350
rect 579498 580294 579554 580350
rect 579622 580294 579678 580350
rect 579250 580170 579306 580226
rect 579374 580170 579430 580226
rect 579498 580170 579554 580226
rect 579622 580170 579678 580226
rect 579250 580046 579306 580102
rect 579374 580046 579430 580102
rect 579498 580046 579554 580102
rect 579622 580046 579678 580102
rect 579250 579922 579306 579978
rect 579374 579922 579430 579978
rect 579498 579922 579554 579978
rect 579622 579922 579678 579978
rect 579250 562294 579306 562350
rect 579374 562294 579430 562350
rect 579498 562294 579554 562350
rect 579622 562294 579678 562350
rect 579250 562170 579306 562226
rect 579374 562170 579430 562226
rect 579498 562170 579554 562226
rect 579622 562170 579678 562226
rect 579250 562046 579306 562102
rect 579374 562046 579430 562102
rect 579498 562046 579554 562102
rect 579622 562046 579678 562102
rect 579250 561922 579306 561978
rect 579374 561922 579430 561978
rect 579498 561922 579554 561978
rect 579622 561922 579678 561978
rect 579250 544294 579306 544350
rect 579374 544294 579430 544350
rect 579498 544294 579554 544350
rect 579622 544294 579678 544350
rect 579250 544170 579306 544226
rect 579374 544170 579430 544226
rect 579498 544170 579554 544226
rect 579622 544170 579678 544226
rect 579250 544046 579306 544102
rect 579374 544046 579430 544102
rect 579498 544046 579554 544102
rect 579622 544046 579678 544102
rect 579250 543922 579306 543978
rect 579374 543922 579430 543978
rect 579498 543922 579554 543978
rect 579622 543922 579678 543978
rect 579250 526294 579306 526350
rect 579374 526294 579430 526350
rect 579498 526294 579554 526350
rect 579622 526294 579678 526350
rect 579250 526170 579306 526226
rect 579374 526170 579430 526226
rect 579498 526170 579554 526226
rect 579622 526170 579678 526226
rect 579250 526046 579306 526102
rect 579374 526046 579430 526102
rect 579498 526046 579554 526102
rect 579622 526046 579678 526102
rect 579250 525922 579306 525978
rect 579374 525922 579430 525978
rect 579498 525922 579554 525978
rect 579622 525922 579678 525978
rect 579250 508294 579306 508350
rect 579374 508294 579430 508350
rect 579498 508294 579554 508350
rect 579622 508294 579678 508350
rect 579250 508170 579306 508226
rect 579374 508170 579430 508226
rect 579498 508170 579554 508226
rect 579622 508170 579678 508226
rect 579250 508046 579306 508102
rect 579374 508046 579430 508102
rect 579498 508046 579554 508102
rect 579622 508046 579678 508102
rect 579250 507922 579306 507978
rect 579374 507922 579430 507978
rect 579498 507922 579554 507978
rect 579622 507922 579678 507978
rect 579250 490294 579306 490350
rect 579374 490294 579430 490350
rect 579498 490294 579554 490350
rect 579622 490294 579678 490350
rect 579250 490170 579306 490226
rect 579374 490170 579430 490226
rect 579498 490170 579554 490226
rect 579622 490170 579678 490226
rect 579250 490046 579306 490102
rect 579374 490046 579430 490102
rect 579498 490046 579554 490102
rect 579622 490046 579678 490102
rect 579250 489922 579306 489978
rect 579374 489922 579430 489978
rect 579498 489922 579554 489978
rect 579622 489922 579678 489978
rect 579250 472294 579306 472350
rect 579374 472294 579430 472350
rect 579498 472294 579554 472350
rect 579622 472294 579678 472350
rect 579250 472170 579306 472226
rect 579374 472170 579430 472226
rect 579498 472170 579554 472226
rect 579622 472170 579678 472226
rect 579250 472046 579306 472102
rect 579374 472046 579430 472102
rect 579498 472046 579554 472102
rect 579622 472046 579678 472102
rect 579250 471922 579306 471978
rect 579374 471922 579430 471978
rect 579498 471922 579554 471978
rect 579622 471922 579678 471978
rect 579250 454294 579306 454350
rect 579374 454294 579430 454350
rect 579498 454294 579554 454350
rect 579622 454294 579678 454350
rect 579250 454170 579306 454226
rect 579374 454170 579430 454226
rect 579498 454170 579554 454226
rect 579622 454170 579678 454226
rect 579250 454046 579306 454102
rect 579374 454046 579430 454102
rect 579498 454046 579554 454102
rect 579622 454046 579678 454102
rect 579250 453922 579306 453978
rect 579374 453922 579430 453978
rect 579498 453922 579554 453978
rect 579622 453922 579678 453978
rect 579250 436294 579306 436350
rect 579374 436294 579430 436350
rect 579498 436294 579554 436350
rect 579622 436294 579678 436350
rect 579250 436170 579306 436226
rect 579374 436170 579430 436226
rect 579498 436170 579554 436226
rect 579622 436170 579678 436226
rect 579250 436046 579306 436102
rect 579374 436046 579430 436102
rect 579498 436046 579554 436102
rect 579622 436046 579678 436102
rect 579250 435922 579306 435978
rect 579374 435922 579430 435978
rect 579498 435922 579554 435978
rect 579622 435922 579678 435978
rect 579250 418294 579306 418350
rect 579374 418294 579430 418350
rect 579498 418294 579554 418350
rect 579622 418294 579678 418350
rect 579250 418170 579306 418226
rect 579374 418170 579430 418226
rect 579498 418170 579554 418226
rect 579622 418170 579678 418226
rect 579250 418046 579306 418102
rect 579374 418046 579430 418102
rect 579498 418046 579554 418102
rect 579622 418046 579678 418102
rect 579250 417922 579306 417978
rect 579374 417922 579430 417978
rect 579498 417922 579554 417978
rect 579622 417922 579678 417978
rect 579250 400294 579306 400350
rect 579374 400294 579430 400350
rect 579498 400294 579554 400350
rect 579622 400294 579678 400350
rect 579250 400170 579306 400226
rect 579374 400170 579430 400226
rect 579498 400170 579554 400226
rect 579622 400170 579678 400226
rect 579250 400046 579306 400102
rect 579374 400046 579430 400102
rect 579498 400046 579554 400102
rect 579622 400046 579678 400102
rect 579250 399922 579306 399978
rect 579374 399922 579430 399978
rect 579498 399922 579554 399978
rect 579622 399922 579678 399978
rect 579250 382294 579306 382350
rect 579374 382294 579430 382350
rect 579498 382294 579554 382350
rect 579622 382294 579678 382350
rect 579250 382170 579306 382226
rect 579374 382170 579430 382226
rect 579498 382170 579554 382226
rect 579622 382170 579678 382226
rect 579250 382046 579306 382102
rect 579374 382046 579430 382102
rect 579498 382046 579554 382102
rect 579622 382046 579678 382102
rect 579250 381922 579306 381978
rect 579374 381922 579430 381978
rect 579498 381922 579554 381978
rect 579622 381922 579678 381978
rect 579250 364294 579306 364350
rect 579374 364294 579430 364350
rect 579498 364294 579554 364350
rect 579622 364294 579678 364350
rect 579250 364170 579306 364226
rect 579374 364170 579430 364226
rect 579498 364170 579554 364226
rect 579622 364170 579678 364226
rect 579250 364046 579306 364102
rect 579374 364046 579430 364102
rect 579498 364046 579554 364102
rect 579622 364046 579678 364102
rect 579250 363922 579306 363978
rect 579374 363922 579430 363978
rect 579498 363922 579554 363978
rect 579622 363922 579678 363978
rect 579250 346294 579306 346350
rect 579374 346294 579430 346350
rect 579498 346294 579554 346350
rect 579622 346294 579678 346350
rect 579250 346170 579306 346226
rect 579374 346170 579430 346226
rect 579498 346170 579554 346226
rect 579622 346170 579678 346226
rect 579250 346046 579306 346102
rect 579374 346046 579430 346102
rect 579498 346046 579554 346102
rect 579622 346046 579678 346102
rect 579250 345922 579306 345978
rect 579374 345922 579430 345978
rect 579498 345922 579554 345978
rect 579622 345922 579678 345978
rect 579250 328294 579306 328350
rect 579374 328294 579430 328350
rect 579498 328294 579554 328350
rect 579622 328294 579678 328350
rect 579250 328170 579306 328226
rect 579374 328170 579430 328226
rect 579498 328170 579554 328226
rect 579622 328170 579678 328226
rect 579250 328046 579306 328102
rect 579374 328046 579430 328102
rect 579498 328046 579554 328102
rect 579622 328046 579678 328102
rect 579250 327922 579306 327978
rect 579374 327922 579430 327978
rect 579498 327922 579554 327978
rect 579622 327922 579678 327978
rect 579250 310294 579306 310350
rect 579374 310294 579430 310350
rect 579498 310294 579554 310350
rect 579622 310294 579678 310350
rect 579250 310170 579306 310226
rect 579374 310170 579430 310226
rect 579498 310170 579554 310226
rect 579622 310170 579678 310226
rect 579250 310046 579306 310102
rect 579374 310046 579430 310102
rect 579498 310046 579554 310102
rect 579622 310046 579678 310102
rect 579250 309922 579306 309978
rect 579374 309922 579430 309978
rect 579498 309922 579554 309978
rect 579622 309922 579678 309978
rect 579250 292294 579306 292350
rect 579374 292294 579430 292350
rect 579498 292294 579554 292350
rect 579622 292294 579678 292350
rect 579250 292170 579306 292226
rect 579374 292170 579430 292226
rect 579498 292170 579554 292226
rect 579622 292170 579678 292226
rect 579250 292046 579306 292102
rect 579374 292046 579430 292102
rect 579498 292046 579554 292102
rect 579622 292046 579678 292102
rect 579250 291922 579306 291978
rect 579374 291922 579430 291978
rect 579498 291922 579554 291978
rect 579622 291922 579678 291978
rect 579250 274294 579306 274350
rect 579374 274294 579430 274350
rect 579498 274294 579554 274350
rect 579622 274294 579678 274350
rect 579250 274170 579306 274226
rect 579374 274170 579430 274226
rect 579498 274170 579554 274226
rect 579622 274170 579678 274226
rect 579250 274046 579306 274102
rect 579374 274046 579430 274102
rect 579498 274046 579554 274102
rect 579622 274046 579678 274102
rect 579250 273922 579306 273978
rect 579374 273922 579430 273978
rect 579498 273922 579554 273978
rect 579622 273922 579678 273978
rect 579250 256294 579306 256350
rect 579374 256294 579430 256350
rect 579498 256294 579554 256350
rect 579622 256294 579678 256350
rect 579250 256170 579306 256226
rect 579374 256170 579430 256226
rect 579498 256170 579554 256226
rect 579622 256170 579678 256226
rect 579250 256046 579306 256102
rect 579374 256046 579430 256102
rect 579498 256046 579554 256102
rect 579622 256046 579678 256102
rect 579250 255922 579306 255978
rect 579374 255922 579430 255978
rect 579498 255922 579554 255978
rect 579622 255922 579678 255978
rect 579250 238294 579306 238350
rect 579374 238294 579430 238350
rect 579498 238294 579554 238350
rect 579622 238294 579678 238350
rect 579250 238170 579306 238226
rect 579374 238170 579430 238226
rect 579498 238170 579554 238226
rect 579622 238170 579678 238226
rect 579250 238046 579306 238102
rect 579374 238046 579430 238102
rect 579498 238046 579554 238102
rect 579622 238046 579678 238102
rect 579250 237922 579306 237978
rect 579374 237922 579430 237978
rect 579498 237922 579554 237978
rect 579622 237922 579678 237978
rect 579250 220294 579306 220350
rect 579374 220294 579430 220350
rect 579498 220294 579554 220350
rect 579622 220294 579678 220350
rect 579250 220170 579306 220226
rect 579374 220170 579430 220226
rect 579498 220170 579554 220226
rect 579622 220170 579678 220226
rect 579250 220046 579306 220102
rect 579374 220046 579430 220102
rect 579498 220046 579554 220102
rect 579622 220046 579678 220102
rect 579250 219922 579306 219978
rect 579374 219922 579430 219978
rect 579498 219922 579554 219978
rect 579622 219922 579678 219978
rect 579250 202294 579306 202350
rect 579374 202294 579430 202350
rect 579498 202294 579554 202350
rect 579622 202294 579678 202350
rect 579250 202170 579306 202226
rect 579374 202170 579430 202226
rect 579498 202170 579554 202226
rect 579622 202170 579678 202226
rect 579250 202046 579306 202102
rect 579374 202046 579430 202102
rect 579498 202046 579554 202102
rect 579622 202046 579678 202102
rect 579250 201922 579306 201978
rect 579374 201922 579430 201978
rect 579498 201922 579554 201978
rect 579622 201922 579678 201978
rect 579250 184294 579306 184350
rect 579374 184294 579430 184350
rect 579498 184294 579554 184350
rect 579622 184294 579678 184350
rect 579250 184170 579306 184226
rect 579374 184170 579430 184226
rect 579498 184170 579554 184226
rect 579622 184170 579678 184226
rect 579250 184046 579306 184102
rect 579374 184046 579430 184102
rect 579498 184046 579554 184102
rect 579622 184046 579678 184102
rect 579250 183922 579306 183978
rect 579374 183922 579430 183978
rect 579498 183922 579554 183978
rect 579622 183922 579678 183978
rect 579250 166294 579306 166350
rect 579374 166294 579430 166350
rect 579498 166294 579554 166350
rect 579622 166294 579678 166350
rect 579250 166170 579306 166226
rect 579374 166170 579430 166226
rect 579498 166170 579554 166226
rect 579622 166170 579678 166226
rect 579250 166046 579306 166102
rect 579374 166046 579430 166102
rect 579498 166046 579554 166102
rect 579622 166046 579678 166102
rect 579250 165922 579306 165978
rect 579374 165922 579430 165978
rect 579498 165922 579554 165978
rect 579622 165922 579678 165978
rect 579250 148294 579306 148350
rect 579374 148294 579430 148350
rect 579498 148294 579554 148350
rect 579622 148294 579678 148350
rect 579250 148170 579306 148226
rect 579374 148170 579430 148226
rect 579498 148170 579554 148226
rect 579622 148170 579678 148226
rect 579250 148046 579306 148102
rect 579374 148046 579430 148102
rect 579498 148046 579554 148102
rect 579622 148046 579678 148102
rect 579250 147922 579306 147978
rect 579374 147922 579430 147978
rect 579498 147922 579554 147978
rect 579622 147922 579678 147978
rect 579250 130294 579306 130350
rect 579374 130294 579430 130350
rect 579498 130294 579554 130350
rect 579622 130294 579678 130350
rect 579250 130170 579306 130226
rect 579374 130170 579430 130226
rect 579498 130170 579554 130226
rect 579622 130170 579678 130226
rect 579250 130046 579306 130102
rect 579374 130046 579430 130102
rect 579498 130046 579554 130102
rect 579622 130046 579678 130102
rect 579250 129922 579306 129978
rect 579374 129922 579430 129978
rect 579498 129922 579554 129978
rect 579622 129922 579678 129978
rect 579250 112294 579306 112350
rect 579374 112294 579430 112350
rect 579498 112294 579554 112350
rect 579622 112294 579678 112350
rect 579250 112170 579306 112226
rect 579374 112170 579430 112226
rect 579498 112170 579554 112226
rect 579622 112170 579678 112226
rect 579250 112046 579306 112102
rect 579374 112046 579430 112102
rect 579498 112046 579554 112102
rect 579622 112046 579678 112102
rect 579250 111922 579306 111978
rect 579374 111922 579430 111978
rect 579498 111922 579554 111978
rect 579622 111922 579678 111978
rect 579250 94294 579306 94350
rect 579374 94294 579430 94350
rect 579498 94294 579554 94350
rect 579622 94294 579678 94350
rect 579250 94170 579306 94226
rect 579374 94170 579430 94226
rect 579498 94170 579554 94226
rect 579622 94170 579678 94226
rect 579250 94046 579306 94102
rect 579374 94046 579430 94102
rect 579498 94046 579554 94102
rect 579622 94046 579678 94102
rect 579250 93922 579306 93978
rect 579374 93922 579430 93978
rect 579498 93922 579554 93978
rect 579622 93922 579678 93978
rect 579250 76294 579306 76350
rect 579374 76294 579430 76350
rect 579498 76294 579554 76350
rect 579622 76294 579678 76350
rect 579250 76170 579306 76226
rect 579374 76170 579430 76226
rect 579498 76170 579554 76226
rect 579622 76170 579678 76226
rect 579250 76046 579306 76102
rect 579374 76046 579430 76102
rect 579498 76046 579554 76102
rect 579622 76046 579678 76102
rect 579250 75922 579306 75978
rect 579374 75922 579430 75978
rect 579498 75922 579554 75978
rect 579622 75922 579678 75978
rect 579250 58294 579306 58350
rect 579374 58294 579430 58350
rect 579498 58294 579554 58350
rect 579622 58294 579678 58350
rect 579250 58170 579306 58226
rect 579374 58170 579430 58226
rect 579498 58170 579554 58226
rect 579622 58170 579678 58226
rect 579250 58046 579306 58102
rect 579374 58046 579430 58102
rect 579498 58046 579554 58102
rect 579622 58046 579678 58102
rect 579250 57922 579306 57978
rect 579374 57922 579430 57978
rect 579498 57922 579554 57978
rect 579622 57922 579678 57978
rect 579250 40294 579306 40350
rect 579374 40294 579430 40350
rect 579498 40294 579554 40350
rect 579622 40294 579678 40350
rect 579250 40170 579306 40226
rect 579374 40170 579430 40226
rect 579498 40170 579554 40226
rect 579622 40170 579678 40226
rect 579250 40046 579306 40102
rect 579374 40046 579430 40102
rect 579498 40046 579554 40102
rect 579622 40046 579678 40102
rect 579250 39922 579306 39978
rect 579374 39922 579430 39978
rect 579498 39922 579554 39978
rect 579622 39922 579678 39978
rect 579250 22294 579306 22350
rect 579374 22294 579430 22350
rect 579498 22294 579554 22350
rect 579622 22294 579678 22350
rect 579250 22170 579306 22226
rect 579374 22170 579430 22226
rect 579498 22170 579554 22226
rect 579622 22170 579678 22226
rect 579250 22046 579306 22102
rect 579374 22046 579430 22102
rect 579498 22046 579554 22102
rect 579622 22046 579678 22102
rect 579250 21922 579306 21978
rect 579374 21922 579430 21978
rect 579498 21922 579554 21978
rect 579622 21922 579678 21978
rect 579250 4294 579306 4350
rect 579374 4294 579430 4350
rect 579498 4294 579554 4350
rect 579622 4294 579678 4350
rect 579250 4170 579306 4226
rect 579374 4170 579430 4226
rect 579498 4170 579554 4226
rect 579622 4170 579678 4226
rect 579250 4046 579306 4102
rect 579374 4046 579430 4102
rect 579498 4046 579554 4102
rect 579622 4046 579678 4102
rect 579250 3922 579306 3978
rect 579374 3922 579430 3978
rect 579498 3922 579554 3978
rect 579622 3922 579678 3978
rect 579250 -216 579306 -160
rect 579374 -216 579430 -160
rect 579498 -216 579554 -160
rect 579622 -216 579678 -160
rect 579250 -340 579306 -284
rect 579374 -340 579430 -284
rect 579498 -340 579554 -284
rect 579622 -340 579678 -284
rect 579250 -464 579306 -408
rect 579374 -464 579430 -408
rect 579498 -464 579554 -408
rect 579622 -464 579678 -408
rect 579250 -588 579306 -532
rect 579374 -588 579430 -532
rect 579498 -588 579554 -532
rect 579622 -588 579678 -532
rect 582970 598116 583026 598172
rect 583094 598116 583150 598172
rect 583218 598116 583274 598172
rect 583342 598116 583398 598172
rect 582970 597992 583026 598048
rect 583094 597992 583150 598048
rect 583218 597992 583274 598048
rect 583342 597992 583398 598048
rect 582970 597868 583026 597924
rect 583094 597868 583150 597924
rect 583218 597868 583274 597924
rect 583342 597868 583398 597924
rect 582970 597744 583026 597800
rect 583094 597744 583150 597800
rect 583218 597744 583274 597800
rect 583342 597744 583398 597800
rect 597456 598116 597512 598172
rect 597580 598116 597636 598172
rect 597704 598116 597760 598172
rect 597828 598116 597884 598172
rect 597456 597992 597512 598048
rect 597580 597992 597636 598048
rect 597704 597992 597760 598048
rect 597828 597992 597884 598048
rect 597456 597868 597512 597924
rect 597580 597868 597636 597924
rect 597704 597868 597760 597924
rect 597828 597868 597884 597924
rect 597456 597744 597512 597800
rect 597580 597744 597636 597800
rect 597704 597744 597760 597800
rect 597828 597744 597884 597800
rect 582970 586294 583026 586350
rect 583094 586294 583150 586350
rect 583218 586294 583274 586350
rect 583342 586294 583398 586350
rect 582970 586170 583026 586226
rect 583094 586170 583150 586226
rect 583218 586170 583274 586226
rect 583342 586170 583398 586226
rect 582970 586046 583026 586102
rect 583094 586046 583150 586102
rect 583218 586046 583274 586102
rect 583342 586046 583398 586102
rect 582970 585922 583026 585978
rect 583094 585922 583150 585978
rect 583218 585922 583274 585978
rect 583342 585922 583398 585978
rect 582970 568294 583026 568350
rect 583094 568294 583150 568350
rect 583218 568294 583274 568350
rect 583342 568294 583398 568350
rect 582970 568170 583026 568226
rect 583094 568170 583150 568226
rect 583218 568170 583274 568226
rect 583342 568170 583398 568226
rect 582970 568046 583026 568102
rect 583094 568046 583150 568102
rect 583218 568046 583274 568102
rect 583342 568046 583398 568102
rect 582970 567922 583026 567978
rect 583094 567922 583150 567978
rect 583218 567922 583274 567978
rect 583342 567922 583398 567978
rect 582970 550294 583026 550350
rect 583094 550294 583150 550350
rect 583218 550294 583274 550350
rect 583342 550294 583398 550350
rect 582970 550170 583026 550226
rect 583094 550170 583150 550226
rect 583218 550170 583274 550226
rect 583342 550170 583398 550226
rect 582970 550046 583026 550102
rect 583094 550046 583150 550102
rect 583218 550046 583274 550102
rect 583342 550046 583398 550102
rect 582970 549922 583026 549978
rect 583094 549922 583150 549978
rect 583218 549922 583274 549978
rect 583342 549922 583398 549978
rect 582970 532294 583026 532350
rect 583094 532294 583150 532350
rect 583218 532294 583274 532350
rect 583342 532294 583398 532350
rect 582970 532170 583026 532226
rect 583094 532170 583150 532226
rect 583218 532170 583274 532226
rect 583342 532170 583398 532226
rect 582970 532046 583026 532102
rect 583094 532046 583150 532102
rect 583218 532046 583274 532102
rect 583342 532046 583398 532102
rect 582970 531922 583026 531978
rect 583094 531922 583150 531978
rect 583218 531922 583274 531978
rect 583342 531922 583398 531978
rect 582970 514294 583026 514350
rect 583094 514294 583150 514350
rect 583218 514294 583274 514350
rect 583342 514294 583398 514350
rect 582970 514170 583026 514226
rect 583094 514170 583150 514226
rect 583218 514170 583274 514226
rect 583342 514170 583398 514226
rect 582970 514046 583026 514102
rect 583094 514046 583150 514102
rect 583218 514046 583274 514102
rect 583342 514046 583398 514102
rect 582970 513922 583026 513978
rect 583094 513922 583150 513978
rect 583218 513922 583274 513978
rect 583342 513922 583398 513978
rect 582970 496294 583026 496350
rect 583094 496294 583150 496350
rect 583218 496294 583274 496350
rect 583342 496294 583398 496350
rect 582970 496170 583026 496226
rect 583094 496170 583150 496226
rect 583218 496170 583274 496226
rect 583342 496170 583398 496226
rect 582970 496046 583026 496102
rect 583094 496046 583150 496102
rect 583218 496046 583274 496102
rect 583342 496046 583398 496102
rect 582970 495922 583026 495978
rect 583094 495922 583150 495978
rect 583218 495922 583274 495978
rect 583342 495922 583398 495978
rect 582970 478294 583026 478350
rect 583094 478294 583150 478350
rect 583218 478294 583274 478350
rect 583342 478294 583398 478350
rect 582970 478170 583026 478226
rect 583094 478170 583150 478226
rect 583218 478170 583274 478226
rect 583342 478170 583398 478226
rect 582970 478046 583026 478102
rect 583094 478046 583150 478102
rect 583218 478046 583274 478102
rect 583342 478046 583398 478102
rect 582970 477922 583026 477978
rect 583094 477922 583150 477978
rect 583218 477922 583274 477978
rect 583342 477922 583398 477978
rect 582970 460294 583026 460350
rect 583094 460294 583150 460350
rect 583218 460294 583274 460350
rect 583342 460294 583398 460350
rect 582970 460170 583026 460226
rect 583094 460170 583150 460226
rect 583218 460170 583274 460226
rect 583342 460170 583398 460226
rect 582970 460046 583026 460102
rect 583094 460046 583150 460102
rect 583218 460046 583274 460102
rect 583342 460046 583398 460102
rect 582970 459922 583026 459978
rect 583094 459922 583150 459978
rect 583218 459922 583274 459978
rect 583342 459922 583398 459978
rect 582970 442294 583026 442350
rect 583094 442294 583150 442350
rect 583218 442294 583274 442350
rect 583342 442294 583398 442350
rect 582970 442170 583026 442226
rect 583094 442170 583150 442226
rect 583218 442170 583274 442226
rect 583342 442170 583398 442226
rect 582970 442046 583026 442102
rect 583094 442046 583150 442102
rect 583218 442046 583274 442102
rect 583342 442046 583398 442102
rect 582970 441922 583026 441978
rect 583094 441922 583150 441978
rect 583218 441922 583274 441978
rect 583342 441922 583398 441978
rect 582970 424294 583026 424350
rect 583094 424294 583150 424350
rect 583218 424294 583274 424350
rect 583342 424294 583398 424350
rect 582970 424170 583026 424226
rect 583094 424170 583150 424226
rect 583218 424170 583274 424226
rect 583342 424170 583398 424226
rect 582970 424046 583026 424102
rect 583094 424046 583150 424102
rect 583218 424046 583274 424102
rect 583342 424046 583398 424102
rect 582970 423922 583026 423978
rect 583094 423922 583150 423978
rect 583218 423922 583274 423978
rect 583342 423922 583398 423978
rect 582970 406294 583026 406350
rect 583094 406294 583150 406350
rect 583218 406294 583274 406350
rect 583342 406294 583398 406350
rect 582970 406170 583026 406226
rect 583094 406170 583150 406226
rect 583218 406170 583274 406226
rect 583342 406170 583398 406226
rect 582970 406046 583026 406102
rect 583094 406046 583150 406102
rect 583218 406046 583274 406102
rect 583342 406046 583398 406102
rect 582970 405922 583026 405978
rect 583094 405922 583150 405978
rect 583218 405922 583274 405978
rect 583342 405922 583398 405978
rect 582970 388294 583026 388350
rect 583094 388294 583150 388350
rect 583218 388294 583274 388350
rect 583342 388294 583398 388350
rect 582970 388170 583026 388226
rect 583094 388170 583150 388226
rect 583218 388170 583274 388226
rect 583342 388170 583398 388226
rect 582970 388046 583026 388102
rect 583094 388046 583150 388102
rect 583218 388046 583274 388102
rect 583342 388046 583398 388102
rect 582970 387922 583026 387978
rect 583094 387922 583150 387978
rect 583218 387922 583274 387978
rect 583342 387922 583398 387978
rect 582970 370294 583026 370350
rect 583094 370294 583150 370350
rect 583218 370294 583274 370350
rect 583342 370294 583398 370350
rect 582970 370170 583026 370226
rect 583094 370170 583150 370226
rect 583218 370170 583274 370226
rect 583342 370170 583398 370226
rect 582970 370046 583026 370102
rect 583094 370046 583150 370102
rect 583218 370046 583274 370102
rect 583342 370046 583398 370102
rect 582970 369922 583026 369978
rect 583094 369922 583150 369978
rect 583218 369922 583274 369978
rect 583342 369922 583398 369978
rect 582970 352294 583026 352350
rect 583094 352294 583150 352350
rect 583218 352294 583274 352350
rect 583342 352294 583398 352350
rect 582970 352170 583026 352226
rect 583094 352170 583150 352226
rect 583218 352170 583274 352226
rect 583342 352170 583398 352226
rect 582970 352046 583026 352102
rect 583094 352046 583150 352102
rect 583218 352046 583274 352102
rect 583342 352046 583398 352102
rect 582970 351922 583026 351978
rect 583094 351922 583150 351978
rect 583218 351922 583274 351978
rect 583342 351922 583398 351978
rect 582970 334294 583026 334350
rect 583094 334294 583150 334350
rect 583218 334294 583274 334350
rect 583342 334294 583398 334350
rect 582970 334170 583026 334226
rect 583094 334170 583150 334226
rect 583218 334170 583274 334226
rect 583342 334170 583398 334226
rect 582970 334046 583026 334102
rect 583094 334046 583150 334102
rect 583218 334046 583274 334102
rect 583342 334046 583398 334102
rect 582970 333922 583026 333978
rect 583094 333922 583150 333978
rect 583218 333922 583274 333978
rect 583342 333922 583398 333978
rect 582970 316294 583026 316350
rect 583094 316294 583150 316350
rect 583218 316294 583274 316350
rect 583342 316294 583398 316350
rect 582970 316170 583026 316226
rect 583094 316170 583150 316226
rect 583218 316170 583274 316226
rect 583342 316170 583398 316226
rect 582970 316046 583026 316102
rect 583094 316046 583150 316102
rect 583218 316046 583274 316102
rect 583342 316046 583398 316102
rect 582970 315922 583026 315978
rect 583094 315922 583150 315978
rect 583218 315922 583274 315978
rect 583342 315922 583398 315978
rect 582970 298294 583026 298350
rect 583094 298294 583150 298350
rect 583218 298294 583274 298350
rect 583342 298294 583398 298350
rect 582970 298170 583026 298226
rect 583094 298170 583150 298226
rect 583218 298170 583274 298226
rect 583342 298170 583398 298226
rect 582970 298046 583026 298102
rect 583094 298046 583150 298102
rect 583218 298046 583274 298102
rect 583342 298046 583398 298102
rect 582970 297922 583026 297978
rect 583094 297922 583150 297978
rect 583218 297922 583274 297978
rect 583342 297922 583398 297978
rect 582970 280294 583026 280350
rect 583094 280294 583150 280350
rect 583218 280294 583274 280350
rect 583342 280294 583398 280350
rect 582970 280170 583026 280226
rect 583094 280170 583150 280226
rect 583218 280170 583274 280226
rect 583342 280170 583398 280226
rect 582970 280046 583026 280102
rect 583094 280046 583150 280102
rect 583218 280046 583274 280102
rect 583342 280046 583398 280102
rect 582970 279922 583026 279978
rect 583094 279922 583150 279978
rect 583218 279922 583274 279978
rect 583342 279922 583398 279978
rect 582970 262294 583026 262350
rect 583094 262294 583150 262350
rect 583218 262294 583274 262350
rect 583342 262294 583398 262350
rect 582970 262170 583026 262226
rect 583094 262170 583150 262226
rect 583218 262170 583274 262226
rect 583342 262170 583398 262226
rect 582970 262046 583026 262102
rect 583094 262046 583150 262102
rect 583218 262046 583274 262102
rect 583342 262046 583398 262102
rect 582970 261922 583026 261978
rect 583094 261922 583150 261978
rect 583218 261922 583274 261978
rect 583342 261922 583398 261978
rect 582970 244294 583026 244350
rect 583094 244294 583150 244350
rect 583218 244294 583274 244350
rect 583342 244294 583398 244350
rect 582970 244170 583026 244226
rect 583094 244170 583150 244226
rect 583218 244170 583274 244226
rect 583342 244170 583398 244226
rect 582970 244046 583026 244102
rect 583094 244046 583150 244102
rect 583218 244046 583274 244102
rect 583342 244046 583398 244102
rect 582970 243922 583026 243978
rect 583094 243922 583150 243978
rect 583218 243922 583274 243978
rect 583342 243922 583398 243978
rect 582970 226294 583026 226350
rect 583094 226294 583150 226350
rect 583218 226294 583274 226350
rect 583342 226294 583398 226350
rect 582970 226170 583026 226226
rect 583094 226170 583150 226226
rect 583218 226170 583274 226226
rect 583342 226170 583398 226226
rect 582970 226046 583026 226102
rect 583094 226046 583150 226102
rect 583218 226046 583274 226102
rect 583342 226046 583398 226102
rect 582970 225922 583026 225978
rect 583094 225922 583150 225978
rect 583218 225922 583274 225978
rect 583342 225922 583398 225978
rect 582970 208294 583026 208350
rect 583094 208294 583150 208350
rect 583218 208294 583274 208350
rect 583342 208294 583398 208350
rect 582970 208170 583026 208226
rect 583094 208170 583150 208226
rect 583218 208170 583274 208226
rect 583342 208170 583398 208226
rect 582970 208046 583026 208102
rect 583094 208046 583150 208102
rect 583218 208046 583274 208102
rect 583342 208046 583398 208102
rect 582970 207922 583026 207978
rect 583094 207922 583150 207978
rect 583218 207922 583274 207978
rect 583342 207922 583398 207978
rect 582970 190294 583026 190350
rect 583094 190294 583150 190350
rect 583218 190294 583274 190350
rect 583342 190294 583398 190350
rect 582970 190170 583026 190226
rect 583094 190170 583150 190226
rect 583218 190170 583274 190226
rect 583342 190170 583398 190226
rect 582970 190046 583026 190102
rect 583094 190046 583150 190102
rect 583218 190046 583274 190102
rect 583342 190046 583398 190102
rect 582970 189922 583026 189978
rect 583094 189922 583150 189978
rect 583218 189922 583274 189978
rect 583342 189922 583398 189978
rect 582970 172294 583026 172350
rect 583094 172294 583150 172350
rect 583218 172294 583274 172350
rect 583342 172294 583398 172350
rect 582970 172170 583026 172226
rect 583094 172170 583150 172226
rect 583218 172170 583274 172226
rect 583342 172170 583398 172226
rect 582970 172046 583026 172102
rect 583094 172046 583150 172102
rect 583218 172046 583274 172102
rect 583342 172046 583398 172102
rect 582970 171922 583026 171978
rect 583094 171922 583150 171978
rect 583218 171922 583274 171978
rect 583342 171922 583398 171978
rect 582970 154294 583026 154350
rect 583094 154294 583150 154350
rect 583218 154294 583274 154350
rect 583342 154294 583398 154350
rect 582970 154170 583026 154226
rect 583094 154170 583150 154226
rect 583218 154170 583274 154226
rect 583342 154170 583398 154226
rect 582970 154046 583026 154102
rect 583094 154046 583150 154102
rect 583218 154046 583274 154102
rect 583342 154046 583398 154102
rect 582970 153922 583026 153978
rect 583094 153922 583150 153978
rect 583218 153922 583274 153978
rect 583342 153922 583398 153978
rect 582970 136294 583026 136350
rect 583094 136294 583150 136350
rect 583218 136294 583274 136350
rect 583342 136294 583398 136350
rect 582970 136170 583026 136226
rect 583094 136170 583150 136226
rect 583218 136170 583274 136226
rect 583342 136170 583398 136226
rect 582970 136046 583026 136102
rect 583094 136046 583150 136102
rect 583218 136046 583274 136102
rect 583342 136046 583398 136102
rect 582970 135922 583026 135978
rect 583094 135922 583150 135978
rect 583218 135922 583274 135978
rect 583342 135922 583398 135978
rect 582970 118294 583026 118350
rect 583094 118294 583150 118350
rect 583218 118294 583274 118350
rect 583342 118294 583398 118350
rect 582970 118170 583026 118226
rect 583094 118170 583150 118226
rect 583218 118170 583274 118226
rect 583342 118170 583398 118226
rect 582970 118046 583026 118102
rect 583094 118046 583150 118102
rect 583218 118046 583274 118102
rect 583342 118046 583398 118102
rect 582970 117922 583026 117978
rect 583094 117922 583150 117978
rect 583218 117922 583274 117978
rect 583342 117922 583398 117978
rect 582970 100294 583026 100350
rect 583094 100294 583150 100350
rect 583218 100294 583274 100350
rect 583342 100294 583398 100350
rect 582970 100170 583026 100226
rect 583094 100170 583150 100226
rect 583218 100170 583274 100226
rect 583342 100170 583398 100226
rect 582970 100046 583026 100102
rect 583094 100046 583150 100102
rect 583218 100046 583274 100102
rect 583342 100046 583398 100102
rect 582970 99922 583026 99978
rect 583094 99922 583150 99978
rect 583218 99922 583274 99978
rect 583342 99922 583398 99978
rect 582970 82294 583026 82350
rect 583094 82294 583150 82350
rect 583218 82294 583274 82350
rect 583342 82294 583398 82350
rect 582970 82170 583026 82226
rect 583094 82170 583150 82226
rect 583218 82170 583274 82226
rect 583342 82170 583398 82226
rect 582970 82046 583026 82102
rect 583094 82046 583150 82102
rect 583218 82046 583274 82102
rect 583342 82046 583398 82102
rect 582970 81922 583026 81978
rect 583094 81922 583150 81978
rect 583218 81922 583274 81978
rect 583342 81922 583398 81978
rect 582970 64294 583026 64350
rect 583094 64294 583150 64350
rect 583218 64294 583274 64350
rect 583342 64294 583398 64350
rect 582970 64170 583026 64226
rect 583094 64170 583150 64226
rect 583218 64170 583274 64226
rect 583342 64170 583398 64226
rect 582970 64046 583026 64102
rect 583094 64046 583150 64102
rect 583218 64046 583274 64102
rect 583342 64046 583398 64102
rect 582970 63922 583026 63978
rect 583094 63922 583150 63978
rect 583218 63922 583274 63978
rect 583342 63922 583398 63978
rect 582970 46294 583026 46350
rect 583094 46294 583150 46350
rect 583218 46294 583274 46350
rect 583342 46294 583398 46350
rect 582970 46170 583026 46226
rect 583094 46170 583150 46226
rect 583218 46170 583274 46226
rect 583342 46170 583398 46226
rect 582970 46046 583026 46102
rect 583094 46046 583150 46102
rect 583218 46046 583274 46102
rect 583342 46046 583398 46102
rect 582970 45922 583026 45978
rect 583094 45922 583150 45978
rect 583218 45922 583274 45978
rect 583342 45922 583398 45978
rect 582970 28294 583026 28350
rect 583094 28294 583150 28350
rect 583218 28294 583274 28350
rect 583342 28294 583398 28350
rect 582970 28170 583026 28226
rect 583094 28170 583150 28226
rect 583218 28170 583274 28226
rect 583342 28170 583398 28226
rect 582970 28046 583026 28102
rect 583094 28046 583150 28102
rect 583218 28046 583274 28102
rect 583342 28046 583398 28102
rect 582970 27922 583026 27978
rect 583094 27922 583150 27978
rect 583218 27922 583274 27978
rect 583342 27922 583398 27978
rect 582970 10294 583026 10350
rect 583094 10294 583150 10350
rect 583218 10294 583274 10350
rect 583342 10294 583398 10350
rect 582970 10170 583026 10226
rect 583094 10170 583150 10226
rect 583218 10170 583274 10226
rect 583342 10170 583398 10226
rect 582970 10046 583026 10102
rect 583094 10046 583150 10102
rect 583218 10046 583274 10102
rect 583342 10046 583398 10102
rect 582970 9922 583026 9978
rect 583094 9922 583150 9978
rect 583218 9922 583274 9978
rect 583342 9922 583398 9978
rect 596496 597156 596552 597212
rect 596620 597156 596676 597212
rect 596744 597156 596800 597212
rect 596868 597156 596924 597212
rect 596496 597032 596552 597088
rect 596620 597032 596676 597088
rect 596744 597032 596800 597088
rect 596868 597032 596924 597088
rect 596496 596908 596552 596964
rect 596620 596908 596676 596964
rect 596744 596908 596800 596964
rect 596868 596908 596924 596964
rect 596496 596784 596552 596840
rect 596620 596784 596676 596840
rect 596744 596784 596800 596840
rect 596868 596784 596924 596840
rect 596496 580294 596552 580350
rect 596620 580294 596676 580350
rect 596744 580294 596800 580350
rect 596868 580294 596924 580350
rect 596496 580170 596552 580226
rect 596620 580170 596676 580226
rect 596744 580170 596800 580226
rect 596868 580170 596924 580226
rect 596496 580046 596552 580102
rect 596620 580046 596676 580102
rect 596744 580046 596800 580102
rect 596868 580046 596924 580102
rect 596496 579922 596552 579978
rect 596620 579922 596676 579978
rect 596744 579922 596800 579978
rect 596868 579922 596924 579978
rect 596496 562294 596552 562350
rect 596620 562294 596676 562350
rect 596744 562294 596800 562350
rect 596868 562294 596924 562350
rect 596496 562170 596552 562226
rect 596620 562170 596676 562226
rect 596744 562170 596800 562226
rect 596868 562170 596924 562226
rect 596496 562046 596552 562102
rect 596620 562046 596676 562102
rect 596744 562046 596800 562102
rect 596868 562046 596924 562102
rect 596496 561922 596552 561978
rect 596620 561922 596676 561978
rect 596744 561922 596800 561978
rect 596868 561922 596924 561978
rect 596496 544294 596552 544350
rect 596620 544294 596676 544350
rect 596744 544294 596800 544350
rect 596868 544294 596924 544350
rect 596496 544170 596552 544226
rect 596620 544170 596676 544226
rect 596744 544170 596800 544226
rect 596868 544170 596924 544226
rect 596496 544046 596552 544102
rect 596620 544046 596676 544102
rect 596744 544046 596800 544102
rect 596868 544046 596924 544102
rect 596496 543922 596552 543978
rect 596620 543922 596676 543978
rect 596744 543922 596800 543978
rect 596868 543922 596924 543978
rect 596496 526294 596552 526350
rect 596620 526294 596676 526350
rect 596744 526294 596800 526350
rect 596868 526294 596924 526350
rect 596496 526170 596552 526226
rect 596620 526170 596676 526226
rect 596744 526170 596800 526226
rect 596868 526170 596924 526226
rect 596496 526046 596552 526102
rect 596620 526046 596676 526102
rect 596744 526046 596800 526102
rect 596868 526046 596924 526102
rect 596496 525922 596552 525978
rect 596620 525922 596676 525978
rect 596744 525922 596800 525978
rect 596868 525922 596924 525978
rect 596496 508294 596552 508350
rect 596620 508294 596676 508350
rect 596744 508294 596800 508350
rect 596868 508294 596924 508350
rect 596496 508170 596552 508226
rect 596620 508170 596676 508226
rect 596744 508170 596800 508226
rect 596868 508170 596924 508226
rect 596496 508046 596552 508102
rect 596620 508046 596676 508102
rect 596744 508046 596800 508102
rect 596868 508046 596924 508102
rect 596496 507922 596552 507978
rect 596620 507922 596676 507978
rect 596744 507922 596800 507978
rect 596868 507922 596924 507978
rect 596496 490294 596552 490350
rect 596620 490294 596676 490350
rect 596744 490294 596800 490350
rect 596868 490294 596924 490350
rect 596496 490170 596552 490226
rect 596620 490170 596676 490226
rect 596744 490170 596800 490226
rect 596868 490170 596924 490226
rect 596496 490046 596552 490102
rect 596620 490046 596676 490102
rect 596744 490046 596800 490102
rect 596868 490046 596924 490102
rect 596496 489922 596552 489978
rect 596620 489922 596676 489978
rect 596744 489922 596800 489978
rect 596868 489922 596924 489978
rect 596496 472294 596552 472350
rect 596620 472294 596676 472350
rect 596744 472294 596800 472350
rect 596868 472294 596924 472350
rect 596496 472170 596552 472226
rect 596620 472170 596676 472226
rect 596744 472170 596800 472226
rect 596868 472170 596924 472226
rect 596496 472046 596552 472102
rect 596620 472046 596676 472102
rect 596744 472046 596800 472102
rect 596868 472046 596924 472102
rect 596496 471922 596552 471978
rect 596620 471922 596676 471978
rect 596744 471922 596800 471978
rect 596868 471922 596924 471978
rect 596496 454294 596552 454350
rect 596620 454294 596676 454350
rect 596744 454294 596800 454350
rect 596868 454294 596924 454350
rect 596496 454170 596552 454226
rect 596620 454170 596676 454226
rect 596744 454170 596800 454226
rect 596868 454170 596924 454226
rect 596496 454046 596552 454102
rect 596620 454046 596676 454102
rect 596744 454046 596800 454102
rect 596868 454046 596924 454102
rect 596496 453922 596552 453978
rect 596620 453922 596676 453978
rect 596744 453922 596800 453978
rect 596868 453922 596924 453978
rect 596496 436294 596552 436350
rect 596620 436294 596676 436350
rect 596744 436294 596800 436350
rect 596868 436294 596924 436350
rect 596496 436170 596552 436226
rect 596620 436170 596676 436226
rect 596744 436170 596800 436226
rect 596868 436170 596924 436226
rect 596496 436046 596552 436102
rect 596620 436046 596676 436102
rect 596744 436046 596800 436102
rect 596868 436046 596924 436102
rect 596496 435922 596552 435978
rect 596620 435922 596676 435978
rect 596744 435922 596800 435978
rect 596868 435922 596924 435978
rect 596496 418294 596552 418350
rect 596620 418294 596676 418350
rect 596744 418294 596800 418350
rect 596868 418294 596924 418350
rect 596496 418170 596552 418226
rect 596620 418170 596676 418226
rect 596744 418170 596800 418226
rect 596868 418170 596924 418226
rect 596496 418046 596552 418102
rect 596620 418046 596676 418102
rect 596744 418046 596800 418102
rect 596868 418046 596924 418102
rect 596496 417922 596552 417978
rect 596620 417922 596676 417978
rect 596744 417922 596800 417978
rect 596868 417922 596924 417978
rect 596496 400294 596552 400350
rect 596620 400294 596676 400350
rect 596744 400294 596800 400350
rect 596868 400294 596924 400350
rect 596496 400170 596552 400226
rect 596620 400170 596676 400226
rect 596744 400170 596800 400226
rect 596868 400170 596924 400226
rect 596496 400046 596552 400102
rect 596620 400046 596676 400102
rect 596744 400046 596800 400102
rect 596868 400046 596924 400102
rect 596496 399922 596552 399978
rect 596620 399922 596676 399978
rect 596744 399922 596800 399978
rect 596868 399922 596924 399978
rect 596496 382294 596552 382350
rect 596620 382294 596676 382350
rect 596744 382294 596800 382350
rect 596868 382294 596924 382350
rect 596496 382170 596552 382226
rect 596620 382170 596676 382226
rect 596744 382170 596800 382226
rect 596868 382170 596924 382226
rect 596496 382046 596552 382102
rect 596620 382046 596676 382102
rect 596744 382046 596800 382102
rect 596868 382046 596924 382102
rect 596496 381922 596552 381978
rect 596620 381922 596676 381978
rect 596744 381922 596800 381978
rect 596868 381922 596924 381978
rect 596496 364294 596552 364350
rect 596620 364294 596676 364350
rect 596744 364294 596800 364350
rect 596868 364294 596924 364350
rect 596496 364170 596552 364226
rect 596620 364170 596676 364226
rect 596744 364170 596800 364226
rect 596868 364170 596924 364226
rect 596496 364046 596552 364102
rect 596620 364046 596676 364102
rect 596744 364046 596800 364102
rect 596868 364046 596924 364102
rect 596496 363922 596552 363978
rect 596620 363922 596676 363978
rect 596744 363922 596800 363978
rect 596868 363922 596924 363978
rect 596496 346294 596552 346350
rect 596620 346294 596676 346350
rect 596744 346294 596800 346350
rect 596868 346294 596924 346350
rect 596496 346170 596552 346226
rect 596620 346170 596676 346226
rect 596744 346170 596800 346226
rect 596868 346170 596924 346226
rect 596496 346046 596552 346102
rect 596620 346046 596676 346102
rect 596744 346046 596800 346102
rect 596868 346046 596924 346102
rect 596496 345922 596552 345978
rect 596620 345922 596676 345978
rect 596744 345922 596800 345978
rect 596868 345922 596924 345978
rect 596496 328294 596552 328350
rect 596620 328294 596676 328350
rect 596744 328294 596800 328350
rect 596868 328294 596924 328350
rect 596496 328170 596552 328226
rect 596620 328170 596676 328226
rect 596744 328170 596800 328226
rect 596868 328170 596924 328226
rect 596496 328046 596552 328102
rect 596620 328046 596676 328102
rect 596744 328046 596800 328102
rect 596868 328046 596924 328102
rect 596496 327922 596552 327978
rect 596620 327922 596676 327978
rect 596744 327922 596800 327978
rect 596868 327922 596924 327978
rect 596496 310294 596552 310350
rect 596620 310294 596676 310350
rect 596744 310294 596800 310350
rect 596868 310294 596924 310350
rect 596496 310170 596552 310226
rect 596620 310170 596676 310226
rect 596744 310170 596800 310226
rect 596868 310170 596924 310226
rect 596496 310046 596552 310102
rect 596620 310046 596676 310102
rect 596744 310046 596800 310102
rect 596868 310046 596924 310102
rect 596496 309922 596552 309978
rect 596620 309922 596676 309978
rect 596744 309922 596800 309978
rect 596868 309922 596924 309978
rect 596496 292294 596552 292350
rect 596620 292294 596676 292350
rect 596744 292294 596800 292350
rect 596868 292294 596924 292350
rect 596496 292170 596552 292226
rect 596620 292170 596676 292226
rect 596744 292170 596800 292226
rect 596868 292170 596924 292226
rect 596496 292046 596552 292102
rect 596620 292046 596676 292102
rect 596744 292046 596800 292102
rect 596868 292046 596924 292102
rect 596496 291922 596552 291978
rect 596620 291922 596676 291978
rect 596744 291922 596800 291978
rect 596868 291922 596924 291978
rect 596496 274294 596552 274350
rect 596620 274294 596676 274350
rect 596744 274294 596800 274350
rect 596868 274294 596924 274350
rect 596496 274170 596552 274226
rect 596620 274170 596676 274226
rect 596744 274170 596800 274226
rect 596868 274170 596924 274226
rect 596496 274046 596552 274102
rect 596620 274046 596676 274102
rect 596744 274046 596800 274102
rect 596868 274046 596924 274102
rect 596496 273922 596552 273978
rect 596620 273922 596676 273978
rect 596744 273922 596800 273978
rect 596868 273922 596924 273978
rect 596496 256294 596552 256350
rect 596620 256294 596676 256350
rect 596744 256294 596800 256350
rect 596868 256294 596924 256350
rect 596496 256170 596552 256226
rect 596620 256170 596676 256226
rect 596744 256170 596800 256226
rect 596868 256170 596924 256226
rect 596496 256046 596552 256102
rect 596620 256046 596676 256102
rect 596744 256046 596800 256102
rect 596868 256046 596924 256102
rect 596496 255922 596552 255978
rect 596620 255922 596676 255978
rect 596744 255922 596800 255978
rect 596868 255922 596924 255978
rect 596496 238294 596552 238350
rect 596620 238294 596676 238350
rect 596744 238294 596800 238350
rect 596868 238294 596924 238350
rect 596496 238170 596552 238226
rect 596620 238170 596676 238226
rect 596744 238170 596800 238226
rect 596868 238170 596924 238226
rect 596496 238046 596552 238102
rect 596620 238046 596676 238102
rect 596744 238046 596800 238102
rect 596868 238046 596924 238102
rect 596496 237922 596552 237978
rect 596620 237922 596676 237978
rect 596744 237922 596800 237978
rect 596868 237922 596924 237978
rect 596496 220294 596552 220350
rect 596620 220294 596676 220350
rect 596744 220294 596800 220350
rect 596868 220294 596924 220350
rect 596496 220170 596552 220226
rect 596620 220170 596676 220226
rect 596744 220170 596800 220226
rect 596868 220170 596924 220226
rect 596496 220046 596552 220102
rect 596620 220046 596676 220102
rect 596744 220046 596800 220102
rect 596868 220046 596924 220102
rect 596496 219922 596552 219978
rect 596620 219922 596676 219978
rect 596744 219922 596800 219978
rect 596868 219922 596924 219978
rect 596496 202294 596552 202350
rect 596620 202294 596676 202350
rect 596744 202294 596800 202350
rect 596868 202294 596924 202350
rect 596496 202170 596552 202226
rect 596620 202170 596676 202226
rect 596744 202170 596800 202226
rect 596868 202170 596924 202226
rect 596496 202046 596552 202102
rect 596620 202046 596676 202102
rect 596744 202046 596800 202102
rect 596868 202046 596924 202102
rect 596496 201922 596552 201978
rect 596620 201922 596676 201978
rect 596744 201922 596800 201978
rect 596868 201922 596924 201978
rect 596496 184294 596552 184350
rect 596620 184294 596676 184350
rect 596744 184294 596800 184350
rect 596868 184294 596924 184350
rect 596496 184170 596552 184226
rect 596620 184170 596676 184226
rect 596744 184170 596800 184226
rect 596868 184170 596924 184226
rect 596496 184046 596552 184102
rect 596620 184046 596676 184102
rect 596744 184046 596800 184102
rect 596868 184046 596924 184102
rect 596496 183922 596552 183978
rect 596620 183922 596676 183978
rect 596744 183922 596800 183978
rect 596868 183922 596924 183978
rect 596496 166294 596552 166350
rect 596620 166294 596676 166350
rect 596744 166294 596800 166350
rect 596868 166294 596924 166350
rect 596496 166170 596552 166226
rect 596620 166170 596676 166226
rect 596744 166170 596800 166226
rect 596868 166170 596924 166226
rect 596496 166046 596552 166102
rect 596620 166046 596676 166102
rect 596744 166046 596800 166102
rect 596868 166046 596924 166102
rect 596496 165922 596552 165978
rect 596620 165922 596676 165978
rect 596744 165922 596800 165978
rect 596868 165922 596924 165978
rect 596496 148294 596552 148350
rect 596620 148294 596676 148350
rect 596744 148294 596800 148350
rect 596868 148294 596924 148350
rect 596496 148170 596552 148226
rect 596620 148170 596676 148226
rect 596744 148170 596800 148226
rect 596868 148170 596924 148226
rect 596496 148046 596552 148102
rect 596620 148046 596676 148102
rect 596744 148046 596800 148102
rect 596868 148046 596924 148102
rect 596496 147922 596552 147978
rect 596620 147922 596676 147978
rect 596744 147922 596800 147978
rect 596868 147922 596924 147978
rect 596496 130294 596552 130350
rect 596620 130294 596676 130350
rect 596744 130294 596800 130350
rect 596868 130294 596924 130350
rect 596496 130170 596552 130226
rect 596620 130170 596676 130226
rect 596744 130170 596800 130226
rect 596868 130170 596924 130226
rect 596496 130046 596552 130102
rect 596620 130046 596676 130102
rect 596744 130046 596800 130102
rect 596868 130046 596924 130102
rect 596496 129922 596552 129978
rect 596620 129922 596676 129978
rect 596744 129922 596800 129978
rect 596868 129922 596924 129978
rect 596496 112294 596552 112350
rect 596620 112294 596676 112350
rect 596744 112294 596800 112350
rect 596868 112294 596924 112350
rect 596496 112170 596552 112226
rect 596620 112170 596676 112226
rect 596744 112170 596800 112226
rect 596868 112170 596924 112226
rect 596496 112046 596552 112102
rect 596620 112046 596676 112102
rect 596744 112046 596800 112102
rect 596868 112046 596924 112102
rect 596496 111922 596552 111978
rect 596620 111922 596676 111978
rect 596744 111922 596800 111978
rect 596868 111922 596924 111978
rect 596496 94294 596552 94350
rect 596620 94294 596676 94350
rect 596744 94294 596800 94350
rect 596868 94294 596924 94350
rect 596496 94170 596552 94226
rect 596620 94170 596676 94226
rect 596744 94170 596800 94226
rect 596868 94170 596924 94226
rect 596496 94046 596552 94102
rect 596620 94046 596676 94102
rect 596744 94046 596800 94102
rect 596868 94046 596924 94102
rect 596496 93922 596552 93978
rect 596620 93922 596676 93978
rect 596744 93922 596800 93978
rect 596868 93922 596924 93978
rect 596496 76294 596552 76350
rect 596620 76294 596676 76350
rect 596744 76294 596800 76350
rect 596868 76294 596924 76350
rect 596496 76170 596552 76226
rect 596620 76170 596676 76226
rect 596744 76170 596800 76226
rect 596868 76170 596924 76226
rect 596496 76046 596552 76102
rect 596620 76046 596676 76102
rect 596744 76046 596800 76102
rect 596868 76046 596924 76102
rect 596496 75922 596552 75978
rect 596620 75922 596676 75978
rect 596744 75922 596800 75978
rect 596868 75922 596924 75978
rect 596496 58294 596552 58350
rect 596620 58294 596676 58350
rect 596744 58294 596800 58350
rect 596868 58294 596924 58350
rect 596496 58170 596552 58226
rect 596620 58170 596676 58226
rect 596744 58170 596800 58226
rect 596868 58170 596924 58226
rect 596496 58046 596552 58102
rect 596620 58046 596676 58102
rect 596744 58046 596800 58102
rect 596868 58046 596924 58102
rect 596496 57922 596552 57978
rect 596620 57922 596676 57978
rect 596744 57922 596800 57978
rect 596868 57922 596924 57978
rect 596496 40294 596552 40350
rect 596620 40294 596676 40350
rect 596744 40294 596800 40350
rect 596868 40294 596924 40350
rect 596496 40170 596552 40226
rect 596620 40170 596676 40226
rect 596744 40170 596800 40226
rect 596868 40170 596924 40226
rect 596496 40046 596552 40102
rect 596620 40046 596676 40102
rect 596744 40046 596800 40102
rect 596868 40046 596924 40102
rect 596496 39922 596552 39978
rect 596620 39922 596676 39978
rect 596744 39922 596800 39978
rect 596868 39922 596924 39978
rect 596496 22294 596552 22350
rect 596620 22294 596676 22350
rect 596744 22294 596800 22350
rect 596868 22294 596924 22350
rect 596496 22170 596552 22226
rect 596620 22170 596676 22226
rect 596744 22170 596800 22226
rect 596868 22170 596924 22226
rect 596496 22046 596552 22102
rect 596620 22046 596676 22102
rect 596744 22046 596800 22102
rect 596868 22046 596924 22102
rect 596496 21922 596552 21978
rect 596620 21922 596676 21978
rect 596744 21922 596800 21978
rect 596868 21922 596924 21978
rect 596496 4294 596552 4350
rect 596620 4294 596676 4350
rect 596744 4294 596800 4350
rect 596868 4294 596924 4350
rect 596496 4170 596552 4226
rect 596620 4170 596676 4226
rect 596744 4170 596800 4226
rect 596868 4170 596924 4226
rect 596496 4046 596552 4102
rect 596620 4046 596676 4102
rect 596744 4046 596800 4102
rect 596868 4046 596924 4102
rect 596496 3922 596552 3978
rect 596620 3922 596676 3978
rect 596744 3922 596800 3978
rect 596868 3922 596924 3978
rect 596496 -216 596552 -160
rect 596620 -216 596676 -160
rect 596744 -216 596800 -160
rect 596868 -216 596924 -160
rect 596496 -340 596552 -284
rect 596620 -340 596676 -284
rect 596744 -340 596800 -284
rect 596868 -340 596924 -284
rect 596496 -464 596552 -408
rect 596620 -464 596676 -408
rect 596744 -464 596800 -408
rect 596868 -464 596924 -408
rect 596496 -588 596552 -532
rect 596620 -588 596676 -532
rect 596744 -588 596800 -532
rect 596868 -588 596924 -532
rect 597456 586294 597512 586350
rect 597580 586294 597636 586350
rect 597704 586294 597760 586350
rect 597828 586294 597884 586350
rect 597456 586170 597512 586226
rect 597580 586170 597636 586226
rect 597704 586170 597760 586226
rect 597828 586170 597884 586226
rect 597456 586046 597512 586102
rect 597580 586046 597636 586102
rect 597704 586046 597760 586102
rect 597828 586046 597884 586102
rect 597456 585922 597512 585978
rect 597580 585922 597636 585978
rect 597704 585922 597760 585978
rect 597828 585922 597884 585978
rect 597456 568294 597512 568350
rect 597580 568294 597636 568350
rect 597704 568294 597760 568350
rect 597828 568294 597884 568350
rect 597456 568170 597512 568226
rect 597580 568170 597636 568226
rect 597704 568170 597760 568226
rect 597828 568170 597884 568226
rect 597456 568046 597512 568102
rect 597580 568046 597636 568102
rect 597704 568046 597760 568102
rect 597828 568046 597884 568102
rect 597456 567922 597512 567978
rect 597580 567922 597636 567978
rect 597704 567922 597760 567978
rect 597828 567922 597884 567978
rect 597456 550294 597512 550350
rect 597580 550294 597636 550350
rect 597704 550294 597760 550350
rect 597828 550294 597884 550350
rect 597456 550170 597512 550226
rect 597580 550170 597636 550226
rect 597704 550170 597760 550226
rect 597828 550170 597884 550226
rect 597456 550046 597512 550102
rect 597580 550046 597636 550102
rect 597704 550046 597760 550102
rect 597828 550046 597884 550102
rect 597456 549922 597512 549978
rect 597580 549922 597636 549978
rect 597704 549922 597760 549978
rect 597828 549922 597884 549978
rect 597456 532294 597512 532350
rect 597580 532294 597636 532350
rect 597704 532294 597760 532350
rect 597828 532294 597884 532350
rect 597456 532170 597512 532226
rect 597580 532170 597636 532226
rect 597704 532170 597760 532226
rect 597828 532170 597884 532226
rect 597456 532046 597512 532102
rect 597580 532046 597636 532102
rect 597704 532046 597760 532102
rect 597828 532046 597884 532102
rect 597456 531922 597512 531978
rect 597580 531922 597636 531978
rect 597704 531922 597760 531978
rect 597828 531922 597884 531978
rect 597456 514294 597512 514350
rect 597580 514294 597636 514350
rect 597704 514294 597760 514350
rect 597828 514294 597884 514350
rect 597456 514170 597512 514226
rect 597580 514170 597636 514226
rect 597704 514170 597760 514226
rect 597828 514170 597884 514226
rect 597456 514046 597512 514102
rect 597580 514046 597636 514102
rect 597704 514046 597760 514102
rect 597828 514046 597884 514102
rect 597456 513922 597512 513978
rect 597580 513922 597636 513978
rect 597704 513922 597760 513978
rect 597828 513922 597884 513978
rect 597456 496294 597512 496350
rect 597580 496294 597636 496350
rect 597704 496294 597760 496350
rect 597828 496294 597884 496350
rect 597456 496170 597512 496226
rect 597580 496170 597636 496226
rect 597704 496170 597760 496226
rect 597828 496170 597884 496226
rect 597456 496046 597512 496102
rect 597580 496046 597636 496102
rect 597704 496046 597760 496102
rect 597828 496046 597884 496102
rect 597456 495922 597512 495978
rect 597580 495922 597636 495978
rect 597704 495922 597760 495978
rect 597828 495922 597884 495978
rect 597456 478294 597512 478350
rect 597580 478294 597636 478350
rect 597704 478294 597760 478350
rect 597828 478294 597884 478350
rect 597456 478170 597512 478226
rect 597580 478170 597636 478226
rect 597704 478170 597760 478226
rect 597828 478170 597884 478226
rect 597456 478046 597512 478102
rect 597580 478046 597636 478102
rect 597704 478046 597760 478102
rect 597828 478046 597884 478102
rect 597456 477922 597512 477978
rect 597580 477922 597636 477978
rect 597704 477922 597760 477978
rect 597828 477922 597884 477978
rect 597456 460294 597512 460350
rect 597580 460294 597636 460350
rect 597704 460294 597760 460350
rect 597828 460294 597884 460350
rect 597456 460170 597512 460226
rect 597580 460170 597636 460226
rect 597704 460170 597760 460226
rect 597828 460170 597884 460226
rect 597456 460046 597512 460102
rect 597580 460046 597636 460102
rect 597704 460046 597760 460102
rect 597828 460046 597884 460102
rect 597456 459922 597512 459978
rect 597580 459922 597636 459978
rect 597704 459922 597760 459978
rect 597828 459922 597884 459978
rect 597456 442294 597512 442350
rect 597580 442294 597636 442350
rect 597704 442294 597760 442350
rect 597828 442294 597884 442350
rect 597456 442170 597512 442226
rect 597580 442170 597636 442226
rect 597704 442170 597760 442226
rect 597828 442170 597884 442226
rect 597456 442046 597512 442102
rect 597580 442046 597636 442102
rect 597704 442046 597760 442102
rect 597828 442046 597884 442102
rect 597456 441922 597512 441978
rect 597580 441922 597636 441978
rect 597704 441922 597760 441978
rect 597828 441922 597884 441978
rect 597456 424294 597512 424350
rect 597580 424294 597636 424350
rect 597704 424294 597760 424350
rect 597828 424294 597884 424350
rect 597456 424170 597512 424226
rect 597580 424170 597636 424226
rect 597704 424170 597760 424226
rect 597828 424170 597884 424226
rect 597456 424046 597512 424102
rect 597580 424046 597636 424102
rect 597704 424046 597760 424102
rect 597828 424046 597884 424102
rect 597456 423922 597512 423978
rect 597580 423922 597636 423978
rect 597704 423922 597760 423978
rect 597828 423922 597884 423978
rect 597456 406294 597512 406350
rect 597580 406294 597636 406350
rect 597704 406294 597760 406350
rect 597828 406294 597884 406350
rect 597456 406170 597512 406226
rect 597580 406170 597636 406226
rect 597704 406170 597760 406226
rect 597828 406170 597884 406226
rect 597456 406046 597512 406102
rect 597580 406046 597636 406102
rect 597704 406046 597760 406102
rect 597828 406046 597884 406102
rect 597456 405922 597512 405978
rect 597580 405922 597636 405978
rect 597704 405922 597760 405978
rect 597828 405922 597884 405978
rect 597456 388294 597512 388350
rect 597580 388294 597636 388350
rect 597704 388294 597760 388350
rect 597828 388294 597884 388350
rect 597456 388170 597512 388226
rect 597580 388170 597636 388226
rect 597704 388170 597760 388226
rect 597828 388170 597884 388226
rect 597456 388046 597512 388102
rect 597580 388046 597636 388102
rect 597704 388046 597760 388102
rect 597828 388046 597884 388102
rect 597456 387922 597512 387978
rect 597580 387922 597636 387978
rect 597704 387922 597760 387978
rect 597828 387922 597884 387978
rect 597456 370294 597512 370350
rect 597580 370294 597636 370350
rect 597704 370294 597760 370350
rect 597828 370294 597884 370350
rect 597456 370170 597512 370226
rect 597580 370170 597636 370226
rect 597704 370170 597760 370226
rect 597828 370170 597884 370226
rect 597456 370046 597512 370102
rect 597580 370046 597636 370102
rect 597704 370046 597760 370102
rect 597828 370046 597884 370102
rect 597456 369922 597512 369978
rect 597580 369922 597636 369978
rect 597704 369922 597760 369978
rect 597828 369922 597884 369978
rect 597456 352294 597512 352350
rect 597580 352294 597636 352350
rect 597704 352294 597760 352350
rect 597828 352294 597884 352350
rect 597456 352170 597512 352226
rect 597580 352170 597636 352226
rect 597704 352170 597760 352226
rect 597828 352170 597884 352226
rect 597456 352046 597512 352102
rect 597580 352046 597636 352102
rect 597704 352046 597760 352102
rect 597828 352046 597884 352102
rect 597456 351922 597512 351978
rect 597580 351922 597636 351978
rect 597704 351922 597760 351978
rect 597828 351922 597884 351978
rect 597456 334294 597512 334350
rect 597580 334294 597636 334350
rect 597704 334294 597760 334350
rect 597828 334294 597884 334350
rect 597456 334170 597512 334226
rect 597580 334170 597636 334226
rect 597704 334170 597760 334226
rect 597828 334170 597884 334226
rect 597456 334046 597512 334102
rect 597580 334046 597636 334102
rect 597704 334046 597760 334102
rect 597828 334046 597884 334102
rect 597456 333922 597512 333978
rect 597580 333922 597636 333978
rect 597704 333922 597760 333978
rect 597828 333922 597884 333978
rect 597456 316294 597512 316350
rect 597580 316294 597636 316350
rect 597704 316294 597760 316350
rect 597828 316294 597884 316350
rect 597456 316170 597512 316226
rect 597580 316170 597636 316226
rect 597704 316170 597760 316226
rect 597828 316170 597884 316226
rect 597456 316046 597512 316102
rect 597580 316046 597636 316102
rect 597704 316046 597760 316102
rect 597828 316046 597884 316102
rect 597456 315922 597512 315978
rect 597580 315922 597636 315978
rect 597704 315922 597760 315978
rect 597828 315922 597884 315978
rect 597456 298294 597512 298350
rect 597580 298294 597636 298350
rect 597704 298294 597760 298350
rect 597828 298294 597884 298350
rect 597456 298170 597512 298226
rect 597580 298170 597636 298226
rect 597704 298170 597760 298226
rect 597828 298170 597884 298226
rect 597456 298046 597512 298102
rect 597580 298046 597636 298102
rect 597704 298046 597760 298102
rect 597828 298046 597884 298102
rect 597456 297922 597512 297978
rect 597580 297922 597636 297978
rect 597704 297922 597760 297978
rect 597828 297922 597884 297978
rect 597456 280294 597512 280350
rect 597580 280294 597636 280350
rect 597704 280294 597760 280350
rect 597828 280294 597884 280350
rect 597456 280170 597512 280226
rect 597580 280170 597636 280226
rect 597704 280170 597760 280226
rect 597828 280170 597884 280226
rect 597456 280046 597512 280102
rect 597580 280046 597636 280102
rect 597704 280046 597760 280102
rect 597828 280046 597884 280102
rect 597456 279922 597512 279978
rect 597580 279922 597636 279978
rect 597704 279922 597760 279978
rect 597828 279922 597884 279978
rect 597456 262294 597512 262350
rect 597580 262294 597636 262350
rect 597704 262294 597760 262350
rect 597828 262294 597884 262350
rect 597456 262170 597512 262226
rect 597580 262170 597636 262226
rect 597704 262170 597760 262226
rect 597828 262170 597884 262226
rect 597456 262046 597512 262102
rect 597580 262046 597636 262102
rect 597704 262046 597760 262102
rect 597828 262046 597884 262102
rect 597456 261922 597512 261978
rect 597580 261922 597636 261978
rect 597704 261922 597760 261978
rect 597828 261922 597884 261978
rect 597456 244294 597512 244350
rect 597580 244294 597636 244350
rect 597704 244294 597760 244350
rect 597828 244294 597884 244350
rect 597456 244170 597512 244226
rect 597580 244170 597636 244226
rect 597704 244170 597760 244226
rect 597828 244170 597884 244226
rect 597456 244046 597512 244102
rect 597580 244046 597636 244102
rect 597704 244046 597760 244102
rect 597828 244046 597884 244102
rect 597456 243922 597512 243978
rect 597580 243922 597636 243978
rect 597704 243922 597760 243978
rect 597828 243922 597884 243978
rect 597456 226294 597512 226350
rect 597580 226294 597636 226350
rect 597704 226294 597760 226350
rect 597828 226294 597884 226350
rect 597456 226170 597512 226226
rect 597580 226170 597636 226226
rect 597704 226170 597760 226226
rect 597828 226170 597884 226226
rect 597456 226046 597512 226102
rect 597580 226046 597636 226102
rect 597704 226046 597760 226102
rect 597828 226046 597884 226102
rect 597456 225922 597512 225978
rect 597580 225922 597636 225978
rect 597704 225922 597760 225978
rect 597828 225922 597884 225978
rect 597456 208294 597512 208350
rect 597580 208294 597636 208350
rect 597704 208294 597760 208350
rect 597828 208294 597884 208350
rect 597456 208170 597512 208226
rect 597580 208170 597636 208226
rect 597704 208170 597760 208226
rect 597828 208170 597884 208226
rect 597456 208046 597512 208102
rect 597580 208046 597636 208102
rect 597704 208046 597760 208102
rect 597828 208046 597884 208102
rect 597456 207922 597512 207978
rect 597580 207922 597636 207978
rect 597704 207922 597760 207978
rect 597828 207922 597884 207978
rect 597456 190294 597512 190350
rect 597580 190294 597636 190350
rect 597704 190294 597760 190350
rect 597828 190294 597884 190350
rect 597456 190170 597512 190226
rect 597580 190170 597636 190226
rect 597704 190170 597760 190226
rect 597828 190170 597884 190226
rect 597456 190046 597512 190102
rect 597580 190046 597636 190102
rect 597704 190046 597760 190102
rect 597828 190046 597884 190102
rect 597456 189922 597512 189978
rect 597580 189922 597636 189978
rect 597704 189922 597760 189978
rect 597828 189922 597884 189978
rect 597456 172294 597512 172350
rect 597580 172294 597636 172350
rect 597704 172294 597760 172350
rect 597828 172294 597884 172350
rect 597456 172170 597512 172226
rect 597580 172170 597636 172226
rect 597704 172170 597760 172226
rect 597828 172170 597884 172226
rect 597456 172046 597512 172102
rect 597580 172046 597636 172102
rect 597704 172046 597760 172102
rect 597828 172046 597884 172102
rect 597456 171922 597512 171978
rect 597580 171922 597636 171978
rect 597704 171922 597760 171978
rect 597828 171922 597884 171978
rect 597456 154294 597512 154350
rect 597580 154294 597636 154350
rect 597704 154294 597760 154350
rect 597828 154294 597884 154350
rect 597456 154170 597512 154226
rect 597580 154170 597636 154226
rect 597704 154170 597760 154226
rect 597828 154170 597884 154226
rect 597456 154046 597512 154102
rect 597580 154046 597636 154102
rect 597704 154046 597760 154102
rect 597828 154046 597884 154102
rect 597456 153922 597512 153978
rect 597580 153922 597636 153978
rect 597704 153922 597760 153978
rect 597828 153922 597884 153978
rect 597456 136294 597512 136350
rect 597580 136294 597636 136350
rect 597704 136294 597760 136350
rect 597828 136294 597884 136350
rect 597456 136170 597512 136226
rect 597580 136170 597636 136226
rect 597704 136170 597760 136226
rect 597828 136170 597884 136226
rect 597456 136046 597512 136102
rect 597580 136046 597636 136102
rect 597704 136046 597760 136102
rect 597828 136046 597884 136102
rect 597456 135922 597512 135978
rect 597580 135922 597636 135978
rect 597704 135922 597760 135978
rect 597828 135922 597884 135978
rect 597456 118294 597512 118350
rect 597580 118294 597636 118350
rect 597704 118294 597760 118350
rect 597828 118294 597884 118350
rect 597456 118170 597512 118226
rect 597580 118170 597636 118226
rect 597704 118170 597760 118226
rect 597828 118170 597884 118226
rect 597456 118046 597512 118102
rect 597580 118046 597636 118102
rect 597704 118046 597760 118102
rect 597828 118046 597884 118102
rect 597456 117922 597512 117978
rect 597580 117922 597636 117978
rect 597704 117922 597760 117978
rect 597828 117922 597884 117978
rect 597456 100294 597512 100350
rect 597580 100294 597636 100350
rect 597704 100294 597760 100350
rect 597828 100294 597884 100350
rect 597456 100170 597512 100226
rect 597580 100170 597636 100226
rect 597704 100170 597760 100226
rect 597828 100170 597884 100226
rect 597456 100046 597512 100102
rect 597580 100046 597636 100102
rect 597704 100046 597760 100102
rect 597828 100046 597884 100102
rect 597456 99922 597512 99978
rect 597580 99922 597636 99978
rect 597704 99922 597760 99978
rect 597828 99922 597884 99978
rect 597456 82294 597512 82350
rect 597580 82294 597636 82350
rect 597704 82294 597760 82350
rect 597828 82294 597884 82350
rect 597456 82170 597512 82226
rect 597580 82170 597636 82226
rect 597704 82170 597760 82226
rect 597828 82170 597884 82226
rect 597456 82046 597512 82102
rect 597580 82046 597636 82102
rect 597704 82046 597760 82102
rect 597828 82046 597884 82102
rect 597456 81922 597512 81978
rect 597580 81922 597636 81978
rect 597704 81922 597760 81978
rect 597828 81922 597884 81978
rect 597456 64294 597512 64350
rect 597580 64294 597636 64350
rect 597704 64294 597760 64350
rect 597828 64294 597884 64350
rect 597456 64170 597512 64226
rect 597580 64170 597636 64226
rect 597704 64170 597760 64226
rect 597828 64170 597884 64226
rect 597456 64046 597512 64102
rect 597580 64046 597636 64102
rect 597704 64046 597760 64102
rect 597828 64046 597884 64102
rect 597456 63922 597512 63978
rect 597580 63922 597636 63978
rect 597704 63922 597760 63978
rect 597828 63922 597884 63978
rect 597456 46294 597512 46350
rect 597580 46294 597636 46350
rect 597704 46294 597760 46350
rect 597828 46294 597884 46350
rect 597456 46170 597512 46226
rect 597580 46170 597636 46226
rect 597704 46170 597760 46226
rect 597828 46170 597884 46226
rect 597456 46046 597512 46102
rect 597580 46046 597636 46102
rect 597704 46046 597760 46102
rect 597828 46046 597884 46102
rect 597456 45922 597512 45978
rect 597580 45922 597636 45978
rect 597704 45922 597760 45978
rect 597828 45922 597884 45978
rect 597456 28294 597512 28350
rect 597580 28294 597636 28350
rect 597704 28294 597760 28350
rect 597828 28294 597884 28350
rect 597456 28170 597512 28226
rect 597580 28170 597636 28226
rect 597704 28170 597760 28226
rect 597828 28170 597884 28226
rect 597456 28046 597512 28102
rect 597580 28046 597636 28102
rect 597704 28046 597760 28102
rect 597828 28046 597884 28102
rect 597456 27922 597512 27978
rect 597580 27922 597636 27978
rect 597704 27922 597760 27978
rect 597828 27922 597884 27978
rect 597456 10294 597512 10350
rect 597580 10294 597636 10350
rect 597704 10294 597760 10350
rect 597828 10294 597884 10350
rect 597456 10170 597512 10226
rect 597580 10170 597636 10226
rect 597704 10170 597760 10226
rect 597828 10170 597884 10226
rect 597456 10046 597512 10102
rect 597580 10046 597636 10102
rect 597704 10046 597760 10102
rect 597828 10046 597884 10102
rect 597456 9922 597512 9978
rect 597580 9922 597636 9978
rect 597704 9922 597760 9978
rect 597828 9922 597884 9978
rect 582970 -1176 583026 -1120
rect 583094 -1176 583150 -1120
rect 583218 -1176 583274 -1120
rect 583342 -1176 583398 -1120
rect 582970 -1300 583026 -1244
rect 583094 -1300 583150 -1244
rect 583218 -1300 583274 -1244
rect 583342 -1300 583398 -1244
rect 582970 -1424 583026 -1368
rect 583094 -1424 583150 -1368
rect 583218 -1424 583274 -1368
rect 583342 -1424 583398 -1368
rect 582970 -1548 583026 -1492
rect 583094 -1548 583150 -1492
rect 583218 -1548 583274 -1492
rect 583342 -1548 583398 -1492
rect 597456 -1176 597512 -1120
rect 597580 -1176 597636 -1120
rect 597704 -1176 597760 -1120
rect 597828 -1176 597884 -1120
rect 597456 -1300 597512 -1244
rect 597580 -1300 597636 -1244
rect 597704 -1300 597760 -1244
rect 597828 -1300 597884 -1244
rect 597456 -1424 597512 -1368
rect 597580 -1424 597636 -1368
rect 597704 -1424 597760 -1368
rect 597828 -1424 597884 -1368
rect 597456 -1548 597512 -1492
rect 597580 -1548 597636 -1492
rect 597704 -1548 597760 -1492
rect 597828 -1548 597884 -1492
<< metal5 >>
rect -1916 598172 597980 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 6970 598172
rect 7026 598116 7094 598172
rect 7150 598116 7218 598172
rect 7274 598116 7342 598172
rect 7398 598116 24970 598172
rect 25026 598116 25094 598172
rect 25150 598116 25218 598172
rect 25274 598116 25342 598172
rect 25398 598116 42970 598172
rect 43026 598116 43094 598172
rect 43150 598116 43218 598172
rect 43274 598116 43342 598172
rect 43398 598116 60970 598172
rect 61026 598116 61094 598172
rect 61150 598116 61218 598172
rect 61274 598116 61342 598172
rect 61398 598116 78970 598172
rect 79026 598116 79094 598172
rect 79150 598116 79218 598172
rect 79274 598116 79342 598172
rect 79398 598116 96970 598172
rect 97026 598116 97094 598172
rect 97150 598116 97218 598172
rect 97274 598116 97342 598172
rect 97398 598116 114970 598172
rect 115026 598116 115094 598172
rect 115150 598116 115218 598172
rect 115274 598116 115342 598172
rect 115398 598116 132970 598172
rect 133026 598116 133094 598172
rect 133150 598116 133218 598172
rect 133274 598116 133342 598172
rect 133398 598116 150970 598172
rect 151026 598116 151094 598172
rect 151150 598116 151218 598172
rect 151274 598116 151342 598172
rect 151398 598116 168970 598172
rect 169026 598116 169094 598172
rect 169150 598116 169218 598172
rect 169274 598116 169342 598172
rect 169398 598116 186970 598172
rect 187026 598116 187094 598172
rect 187150 598116 187218 598172
rect 187274 598116 187342 598172
rect 187398 598116 204970 598172
rect 205026 598116 205094 598172
rect 205150 598116 205218 598172
rect 205274 598116 205342 598172
rect 205398 598116 222970 598172
rect 223026 598116 223094 598172
rect 223150 598116 223218 598172
rect 223274 598116 223342 598172
rect 223398 598116 240970 598172
rect 241026 598116 241094 598172
rect 241150 598116 241218 598172
rect 241274 598116 241342 598172
rect 241398 598116 258970 598172
rect 259026 598116 259094 598172
rect 259150 598116 259218 598172
rect 259274 598116 259342 598172
rect 259398 598116 276970 598172
rect 277026 598116 277094 598172
rect 277150 598116 277218 598172
rect 277274 598116 277342 598172
rect 277398 598116 294970 598172
rect 295026 598116 295094 598172
rect 295150 598116 295218 598172
rect 295274 598116 295342 598172
rect 295398 598116 312970 598172
rect 313026 598116 313094 598172
rect 313150 598116 313218 598172
rect 313274 598116 313342 598172
rect 313398 598116 330970 598172
rect 331026 598116 331094 598172
rect 331150 598116 331218 598172
rect 331274 598116 331342 598172
rect 331398 598116 348970 598172
rect 349026 598116 349094 598172
rect 349150 598116 349218 598172
rect 349274 598116 349342 598172
rect 349398 598116 366970 598172
rect 367026 598116 367094 598172
rect 367150 598116 367218 598172
rect 367274 598116 367342 598172
rect 367398 598116 384970 598172
rect 385026 598116 385094 598172
rect 385150 598116 385218 598172
rect 385274 598116 385342 598172
rect 385398 598116 402970 598172
rect 403026 598116 403094 598172
rect 403150 598116 403218 598172
rect 403274 598116 403342 598172
rect 403398 598116 420970 598172
rect 421026 598116 421094 598172
rect 421150 598116 421218 598172
rect 421274 598116 421342 598172
rect 421398 598116 438970 598172
rect 439026 598116 439094 598172
rect 439150 598116 439218 598172
rect 439274 598116 439342 598172
rect 439398 598116 456970 598172
rect 457026 598116 457094 598172
rect 457150 598116 457218 598172
rect 457274 598116 457342 598172
rect 457398 598116 474970 598172
rect 475026 598116 475094 598172
rect 475150 598116 475218 598172
rect 475274 598116 475342 598172
rect 475398 598116 492970 598172
rect 493026 598116 493094 598172
rect 493150 598116 493218 598172
rect 493274 598116 493342 598172
rect 493398 598116 510970 598172
rect 511026 598116 511094 598172
rect 511150 598116 511218 598172
rect 511274 598116 511342 598172
rect 511398 598116 528970 598172
rect 529026 598116 529094 598172
rect 529150 598116 529218 598172
rect 529274 598116 529342 598172
rect 529398 598116 546970 598172
rect 547026 598116 547094 598172
rect 547150 598116 547218 598172
rect 547274 598116 547342 598172
rect 547398 598116 564970 598172
rect 565026 598116 565094 598172
rect 565150 598116 565218 598172
rect 565274 598116 565342 598172
rect 565398 598116 582970 598172
rect 583026 598116 583094 598172
rect 583150 598116 583218 598172
rect 583274 598116 583342 598172
rect 583398 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect -1916 598048 597980 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 6970 598048
rect 7026 597992 7094 598048
rect 7150 597992 7218 598048
rect 7274 597992 7342 598048
rect 7398 597992 24970 598048
rect 25026 597992 25094 598048
rect 25150 597992 25218 598048
rect 25274 597992 25342 598048
rect 25398 597992 42970 598048
rect 43026 597992 43094 598048
rect 43150 597992 43218 598048
rect 43274 597992 43342 598048
rect 43398 597992 60970 598048
rect 61026 597992 61094 598048
rect 61150 597992 61218 598048
rect 61274 597992 61342 598048
rect 61398 597992 78970 598048
rect 79026 597992 79094 598048
rect 79150 597992 79218 598048
rect 79274 597992 79342 598048
rect 79398 597992 96970 598048
rect 97026 597992 97094 598048
rect 97150 597992 97218 598048
rect 97274 597992 97342 598048
rect 97398 597992 114970 598048
rect 115026 597992 115094 598048
rect 115150 597992 115218 598048
rect 115274 597992 115342 598048
rect 115398 597992 132970 598048
rect 133026 597992 133094 598048
rect 133150 597992 133218 598048
rect 133274 597992 133342 598048
rect 133398 597992 150970 598048
rect 151026 597992 151094 598048
rect 151150 597992 151218 598048
rect 151274 597992 151342 598048
rect 151398 597992 168970 598048
rect 169026 597992 169094 598048
rect 169150 597992 169218 598048
rect 169274 597992 169342 598048
rect 169398 597992 186970 598048
rect 187026 597992 187094 598048
rect 187150 597992 187218 598048
rect 187274 597992 187342 598048
rect 187398 597992 204970 598048
rect 205026 597992 205094 598048
rect 205150 597992 205218 598048
rect 205274 597992 205342 598048
rect 205398 597992 222970 598048
rect 223026 597992 223094 598048
rect 223150 597992 223218 598048
rect 223274 597992 223342 598048
rect 223398 597992 240970 598048
rect 241026 597992 241094 598048
rect 241150 597992 241218 598048
rect 241274 597992 241342 598048
rect 241398 597992 258970 598048
rect 259026 597992 259094 598048
rect 259150 597992 259218 598048
rect 259274 597992 259342 598048
rect 259398 597992 276970 598048
rect 277026 597992 277094 598048
rect 277150 597992 277218 598048
rect 277274 597992 277342 598048
rect 277398 597992 294970 598048
rect 295026 597992 295094 598048
rect 295150 597992 295218 598048
rect 295274 597992 295342 598048
rect 295398 597992 312970 598048
rect 313026 597992 313094 598048
rect 313150 597992 313218 598048
rect 313274 597992 313342 598048
rect 313398 597992 330970 598048
rect 331026 597992 331094 598048
rect 331150 597992 331218 598048
rect 331274 597992 331342 598048
rect 331398 597992 348970 598048
rect 349026 597992 349094 598048
rect 349150 597992 349218 598048
rect 349274 597992 349342 598048
rect 349398 597992 366970 598048
rect 367026 597992 367094 598048
rect 367150 597992 367218 598048
rect 367274 597992 367342 598048
rect 367398 597992 384970 598048
rect 385026 597992 385094 598048
rect 385150 597992 385218 598048
rect 385274 597992 385342 598048
rect 385398 597992 402970 598048
rect 403026 597992 403094 598048
rect 403150 597992 403218 598048
rect 403274 597992 403342 598048
rect 403398 597992 420970 598048
rect 421026 597992 421094 598048
rect 421150 597992 421218 598048
rect 421274 597992 421342 598048
rect 421398 597992 438970 598048
rect 439026 597992 439094 598048
rect 439150 597992 439218 598048
rect 439274 597992 439342 598048
rect 439398 597992 456970 598048
rect 457026 597992 457094 598048
rect 457150 597992 457218 598048
rect 457274 597992 457342 598048
rect 457398 597992 474970 598048
rect 475026 597992 475094 598048
rect 475150 597992 475218 598048
rect 475274 597992 475342 598048
rect 475398 597992 492970 598048
rect 493026 597992 493094 598048
rect 493150 597992 493218 598048
rect 493274 597992 493342 598048
rect 493398 597992 510970 598048
rect 511026 597992 511094 598048
rect 511150 597992 511218 598048
rect 511274 597992 511342 598048
rect 511398 597992 528970 598048
rect 529026 597992 529094 598048
rect 529150 597992 529218 598048
rect 529274 597992 529342 598048
rect 529398 597992 546970 598048
rect 547026 597992 547094 598048
rect 547150 597992 547218 598048
rect 547274 597992 547342 598048
rect 547398 597992 564970 598048
rect 565026 597992 565094 598048
rect 565150 597992 565218 598048
rect 565274 597992 565342 598048
rect 565398 597992 582970 598048
rect 583026 597992 583094 598048
rect 583150 597992 583218 598048
rect 583274 597992 583342 598048
rect 583398 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect -1916 597924 597980 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 6970 597924
rect 7026 597868 7094 597924
rect 7150 597868 7218 597924
rect 7274 597868 7342 597924
rect 7398 597868 24970 597924
rect 25026 597868 25094 597924
rect 25150 597868 25218 597924
rect 25274 597868 25342 597924
rect 25398 597868 42970 597924
rect 43026 597868 43094 597924
rect 43150 597868 43218 597924
rect 43274 597868 43342 597924
rect 43398 597868 60970 597924
rect 61026 597868 61094 597924
rect 61150 597868 61218 597924
rect 61274 597868 61342 597924
rect 61398 597868 78970 597924
rect 79026 597868 79094 597924
rect 79150 597868 79218 597924
rect 79274 597868 79342 597924
rect 79398 597868 96970 597924
rect 97026 597868 97094 597924
rect 97150 597868 97218 597924
rect 97274 597868 97342 597924
rect 97398 597868 114970 597924
rect 115026 597868 115094 597924
rect 115150 597868 115218 597924
rect 115274 597868 115342 597924
rect 115398 597868 132970 597924
rect 133026 597868 133094 597924
rect 133150 597868 133218 597924
rect 133274 597868 133342 597924
rect 133398 597868 150970 597924
rect 151026 597868 151094 597924
rect 151150 597868 151218 597924
rect 151274 597868 151342 597924
rect 151398 597868 168970 597924
rect 169026 597868 169094 597924
rect 169150 597868 169218 597924
rect 169274 597868 169342 597924
rect 169398 597868 186970 597924
rect 187026 597868 187094 597924
rect 187150 597868 187218 597924
rect 187274 597868 187342 597924
rect 187398 597868 204970 597924
rect 205026 597868 205094 597924
rect 205150 597868 205218 597924
rect 205274 597868 205342 597924
rect 205398 597868 222970 597924
rect 223026 597868 223094 597924
rect 223150 597868 223218 597924
rect 223274 597868 223342 597924
rect 223398 597868 240970 597924
rect 241026 597868 241094 597924
rect 241150 597868 241218 597924
rect 241274 597868 241342 597924
rect 241398 597868 258970 597924
rect 259026 597868 259094 597924
rect 259150 597868 259218 597924
rect 259274 597868 259342 597924
rect 259398 597868 276970 597924
rect 277026 597868 277094 597924
rect 277150 597868 277218 597924
rect 277274 597868 277342 597924
rect 277398 597868 294970 597924
rect 295026 597868 295094 597924
rect 295150 597868 295218 597924
rect 295274 597868 295342 597924
rect 295398 597868 312970 597924
rect 313026 597868 313094 597924
rect 313150 597868 313218 597924
rect 313274 597868 313342 597924
rect 313398 597868 330970 597924
rect 331026 597868 331094 597924
rect 331150 597868 331218 597924
rect 331274 597868 331342 597924
rect 331398 597868 348970 597924
rect 349026 597868 349094 597924
rect 349150 597868 349218 597924
rect 349274 597868 349342 597924
rect 349398 597868 366970 597924
rect 367026 597868 367094 597924
rect 367150 597868 367218 597924
rect 367274 597868 367342 597924
rect 367398 597868 384970 597924
rect 385026 597868 385094 597924
rect 385150 597868 385218 597924
rect 385274 597868 385342 597924
rect 385398 597868 402970 597924
rect 403026 597868 403094 597924
rect 403150 597868 403218 597924
rect 403274 597868 403342 597924
rect 403398 597868 420970 597924
rect 421026 597868 421094 597924
rect 421150 597868 421218 597924
rect 421274 597868 421342 597924
rect 421398 597868 438970 597924
rect 439026 597868 439094 597924
rect 439150 597868 439218 597924
rect 439274 597868 439342 597924
rect 439398 597868 456970 597924
rect 457026 597868 457094 597924
rect 457150 597868 457218 597924
rect 457274 597868 457342 597924
rect 457398 597868 474970 597924
rect 475026 597868 475094 597924
rect 475150 597868 475218 597924
rect 475274 597868 475342 597924
rect 475398 597868 492970 597924
rect 493026 597868 493094 597924
rect 493150 597868 493218 597924
rect 493274 597868 493342 597924
rect 493398 597868 510970 597924
rect 511026 597868 511094 597924
rect 511150 597868 511218 597924
rect 511274 597868 511342 597924
rect 511398 597868 528970 597924
rect 529026 597868 529094 597924
rect 529150 597868 529218 597924
rect 529274 597868 529342 597924
rect 529398 597868 546970 597924
rect 547026 597868 547094 597924
rect 547150 597868 547218 597924
rect 547274 597868 547342 597924
rect 547398 597868 564970 597924
rect 565026 597868 565094 597924
rect 565150 597868 565218 597924
rect 565274 597868 565342 597924
rect 565398 597868 582970 597924
rect 583026 597868 583094 597924
rect 583150 597868 583218 597924
rect 583274 597868 583342 597924
rect 583398 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect -1916 597800 597980 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 6970 597800
rect 7026 597744 7094 597800
rect 7150 597744 7218 597800
rect 7274 597744 7342 597800
rect 7398 597744 24970 597800
rect 25026 597744 25094 597800
rect 25150 597744 25218 597800
rect 25274 597744 25342 597800
rect 25398 597744 42970 597800
rect 43026 597744 43094 597800
rect 43150 597744 43218 597800
rect 43274 597744 43342 597800
rect 43398 597744 60970 597800
rect 61026 597744 61094 597800
rect 61150 597744 61218 597800
rect 61274 597744 61342 597800
rect 61398 597744 78970 597800
rect 79026 597744 79094 597800
rect 79150 597744 79218 597800
rect 79274 597744 79342 597800
rect 79398 597744 96970 597800
rect 97026 597744 97094 597800
rect 97150 597744 97218 597800
rect 97274 597744 97342 597800
rect 97398 597744 114970 597800
rect 115026 597744 115094 597800
rect 115150 597744 115218 597800
rect 115274 597744 115342 597800
rect 115398 597744 132970 597800
rect 133026 597744 133094 597800
rect 133150 597744 133218 597800
rect 133274 597744 133342 597800
rect 133398 597744 150970 597800
rect 151026 597744 151094 597800
rect 151150 597744 151218 597800
rect 151274 597744 151342 597800
rect 151398 597744 168970 597800
rect 169026 597744 169094 597800
rect 169150 597744 169218 597800
rect 169274 597744 169342 597800
rect 169398 597744 186970 597800
rect 187026 597744 187094 597800
rect 187150 597744 187218 597800
rect 187274 597744 187342 597800
rect 187398 597744 204970 597800
rect 205026 597744 205094 597800
rect 205150 597744 205218 597800
rect 205274 597744 205342 597800
rect 205398 597744 222970 597800
rect 223026 597744 223094 597800
rect 223150 597744 223218 597800
rect 223274 597744 223342 597800
rect 223398 597744 240970 597800
rect 241026 597744 241094 597800
rect 241150 597744 241218 597800
rect 241274 597744 241342 597800
rect 241398 597744 258970 597800
rect 259026 597744 259094 597800
rect 259150 597744 259218 597800
rect 259274 597744 259342 597800
rect 259398 597744 276970 597800
rect 277026 597744 277094 597800
rect 277150 597744 277218 597800
rect 277274 597744 277342 597800
rect 277398 597744 294970 597800
rect 295026 597744 295094 597800
rect 295150 597744 295218 597800
rect 295274 597744 295342 597800
rect 295398 597744 312970 597800
rect 313026 597744 313094 597800
rect 313150 597744 313218 597800
rect 313274 597744 313342 597800
rect 313398 597744 330970 597800
rect 331026 597744 331094 597800
rect 331150 597744 331218 597800
rect 331274 597744 331342 597800
rect 331398 597744 348970 597800
rect 349026 597744 349094 597800
rect 349150 597744 349218 597800
rect 349274 597744 349342 597800
rect 349398 597744 366970 597800
rect 367026 597744 367094 597800
rect 367150 597744 367218 597800
rect 367274 597744 367342 597800
rect 367398 597744 384970 597800
rect 385026 597744 385094 597800
rect 385150 597744 385218 597800
rect 385274 597744 385342 597800
rect 385398 597744 402970 597800
rect 403026 597744 403094 597800
rect 403150 597744 403218 597800
rect 403274 597744 403342 597800
rect 403398 597744 420970 597800
rect 421026 597744 421094 597800
rect 421150 597744 421218 597800
rect 421274 597744 421342 597800
rect 421398 597744 438970 597800
rect 439026 597744 439094 597800
rect 439150 597744 439218 597800
rect 439274 597744 439342 597800
rect 439398 597744 456970 597800
rect 457026 597744 457094 597800
rect 457150 597744 457218 597800
rect 457274 597744 457342 597800
rect 457398 597744 474970 597800
rect 475026 597744 475094 597800
rect 475150 597744 475218 597800
rect 475274 597744 475342 597800
rect 475398 597744 492970 597800
rect 493026 597744 493094 597800
rect 493150 597744 493218 597800
rect 493274 597744 493342 597800
rect 493398 597744 510970 597800
rect 511026 597744 511094 597800
rect 511150 597744 511218 597800
rect 511274 597744 511342 597800
rect 511398 597744 528970 597800
rect 529026 597744 529094 597800
rect 529150 597744 529218 597800
rect 529274 597744 529342 597800
rect 529398 597744 546970 597800
rect 547026 597744 547094 597800
rect 547150 597744 547218 597800
rect 547274 597744 547342 597800
rect 547398 597744 564970 597800
rect 565026 597744 565094 597800
rect 565150 597744 565218 597800
rect 565274 597744 565342 597800
rect 565398 597744 582970 597800
rect 583026 597744 583094 597800
rect 583150 597744 583218 597800
rect 583274 597744 583342 597800
rect 583398 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect -1916 597648 597980 597744
rect -956 597212 597020 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 3250 597212
rect 3306 597156 3374 597212
rect 3430 597156 3498 597212
rect 3554 597156 3622 597212
rect 3678 597156 21250 597212
rect 21306 597156 21374 597212
rect 21430 597156 21498 597212
rect 21554 597156 21622 597212
rect 21678 597156 39250 597212
rect 39306 597156 39374 597212
rect 39430 597156 39498 597212
rect 39554 597156 39622 597212
rect 39678 597156 57250 597212
rect 57306 597156 57374 597212
rect 57430 597156 57498 597212
rect 57554 597156 57622 597212
rect 57678 597156 75250 597212
rect 75306 597156 75374 597212
rect 75430 597156 75498 597212
rect 75554 597156 75622 597212
rect 75678 597156 93250 597212
rect 93306 597156 93374 597212
rect 93430 597156 93498 597212
rect 93554 597156 93622 597212
rect 93678 597156 111250 597212
rect 111306 597156 111374 597212
rect 111430 597156 111498 597212
rect 111554 597156 111622 597212
rect 111678 597156 129250 597212
rect 129306 597156 129374 597212
rect 129430 597156 129498 597212
rect 129554 597156 129622 597212
rect 129678 597156 147250 597212
rect 147306 597156 147374 597212
rect 147430 597156 147498 597212
rect 147554 597156 147622 597212
rect 147678 597156 165250 597212
rect 165306 597156 165374 597212
rect 165430 597156 165498 597212
rect 165554 597156 165622 597212
rect 165678 597156 183250 597212
rect 183306 597156 183374 597212
rect 183430 597156 183498 597212
rect 183554 597156 183622 597212
rect 183678 597156 201250 597212
rect 201306 597156 201374 597212
rect 201430 597156 201498 597212
rect 201554 597156 201622 597212
rect 201678 597156 219250 597212
rect 219306 597156 219374 597212
rect 219430 597156 219498 597212
rect 219554 597156 219622 597212
rect 219678 597156 237250 597212
rect 237306 597156 237374 597212
rect 237430 597156 237498 597212
rect 237554 597156 237622 597212
rect 237678 597156 255250 597212
rect 255306 597156 255374 597212
rect 255430 597156 255498 597212
rect 255554 597156 255622 597212
rect 255678 597156 273250 597212
rect 273306 597156 273374 597212
rect 273430 597156 273498 597212
rect 273554 597156 273622 597212
rect 273678 597156 291250 597212
rect 291306 597156 291374 597212
rect 291430 597156 291498 597212
rect 291554 597156 291622 597212
rect 291678 597156 309250 597212
rect 309306 597156 309374 597212
rect 309430 597156 309498 597212
rect 309554 597156 309622 597212
rect 309678 597156 327250 597212
rect 327306 597156 327374 597212
rect 327430 597156 327498 597212
rect 327554 597156 327622 597212
rect 327678 597156 345250 597212
rect 345306 597156 345374 597212
rect 345430 597156 345498 597212
rect 345554 597156 345622 597212
rect 345678 597156 363250 597212
rect 363306 597156 363374 597212
rect 363430 597156 363498 597212
rect 363554 597156 363622 597212
rect 363678 597156 381250 597212
rect 381306 597156 381374 597212
rect 381430 597156 381498 597212
rect 381554 597156 381622 597212
rect 381678 597156 399250 597212
rect 399306 597156 399374 597212
rect 399430 597156 399498 597212
rect 399554 597156 399622 597212
rect 399678 597156 417250 597212
rect 417306 597156 417374 597212
rect 417430 597156 417498 597212
rect 417554 597156 417622 597212
rect 417678 597156 435250 597212
rect 435306 597156 435374 597212
rect 435430 597156 435498 597212
rect 435554 597156 435622 597212
rect 435678 597156 453250 597212
rect 453306 597156 453374 597212
rect 453430 597156 453498 597212
rect 453554 597156 453622 597212
rect 453678 597156 471250 597212
rect 471306 597156 471374 597212
rect 471430 597156 471498 597212
rect 471554 597156 471622 597212
rect 471678 597156 489250 597212
rect 489306 597156 489374 597212
rect 489430 597156 489498 597212
rect 489554 597156 489622 597212
rect 489678 597156 507250 597212
rect 507306 597156 507374 597212
rect 507430 597156 507498 597212
rect 507554 597156 507622 597212
rect 507678 597156 525250 597212
rect 525306 597156 525374 597212
rect 525430 597156 525498 597212
rect 525554 597156 525622 597212
rect 525678 597156 543250 597212
rect 543306 597156 543374 597212
rect 543430 597156 543498 597212
rect 543554 597156 543622 597212
rect 543678 597156 561250 597212
rect 561306 597156 561374 597212
rect 561430 597156 561498 597212
rect 561554 597156 561622 597212
rect 561678 597156 579250 597212
rect 579306 597156 579374 597212
rect 579430 597156 579498 597212
rect 579554 597156 579622 597212
rect 579678 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect -956 597088 597020 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 3250 597088
rect 3306 597032 3374 597088
rect 3430 597032 3498 597088
rect 3554 597032 3622 597088
rect 3678 597032 21250 597088
rect 21306 597032 21374 597088
rect 21430 597032 21498 597088
rect 21554 597032 21622 597088
rect 21678 597032 39250 597088
rect 39306 597032 39374 597088
rect 39430 597032 39498 597088
rect 39554 597032 39622 597088
rect 39678 597032 57250 597088
rect 57306 597032 57374 597088
rect 57430 597032 57498 597088
rect 57554 597032 57622 597088
rect 57678 597032 75250 597088
rect 75306 597032 75374 597088
rect 75430 597032 75498 597088
rect 75554 597032 75622 597088
rect 75678 597032 93250 597088
rect 93306 597032 93374 597088
rect 93430 597032 93498 597088
rect 93554 597032 93622 597088
rect 93678 597032 111250 597088
rect 111306 597032 111374 597088
rect 111430 597032 111498 597088
rect 111554 597032 111622 597088
rect 111678 597032 129250 597088
rect 129306 597032 129374 597088
rect 129430 597032 129498 597088
rect 129554 597032 129622 597088
rect 129678 597032 147250 597088
rect 147306 597032 147374 597088
rect 147430 597032 147498 597088
rect 147554 597032 147622 597088
rect 147678 597032 165250 597088
rect 165306 597032 165374 597088
rect 165430 597032 165498 597088
rect 165554 597032 165622 597088
rect 165678 597032 183250 597088
rect 183306 597032 183374 597088
rect 183430 597032 183498 597088
rect 183554 597032 183622 597088
rect 183678 597032 201250 597088
rect 201306 597032 201374 597088
rect 201430 597032 201498 597088
rect 201554 597032 201622 597088
rect 201678 597032 219250 597088
rect 219306 597032 219374 597088
rect 219430 597032 219498 597088
rect 219554 597032 219622 597088
rect 219678 597032 237250 597088
rect 237306 597032 237374 597088
rect 237430 597032 237498 597088
rect 237554 597032 237622 597088
rect 237678 597032 255250 597088
rect 255306 597032 255374 597088
rect 255430 597032 255498 597088
rect 255554 597032 255622 597088
rect 255678 597032 273250 597088
rect 273306 597032 273374 597088
rect 273430 597032 273498 597088
rect 273554 597032 273622 597088
rect 273678 597032 291250 597088
rect 291306 597032 291374 597088
rect 291430 597032 291498 597088
rect 291554 597032 291622 597088
rect 291678 597032 309250 597088
rect 309306 597032 309374 597088
rect 309430 597032 309498 597088
rect 309554 597032 309622 597088
rect 309678 597032 327250 597088
rect 327306 597032 327374 597088
rect 327430 597032 327498 597088
rect 327554 597032 327622 597088
rect 327678 597032 345250 597088
rect 345306 597032 345374 597088
rect 345430 597032 345498 597088
rect 345554 597032 345622 597088
rect 345678 597032 363250 597088
rect 363306 597032 363374 597088
rect 363430 597032 363498 597088
rect 363554 597032 363622 597088
rect 363678 597032 381250 597088
rect 381306 597032 381374 597088
rect 381430 597032 381498 597088
rect 381554 597032 381622 597088
rect 381678 597032 399250 597088
rect 399306 597032 399374 597088
rect 399430 597032 399498 597088
rect 399554 597032 399622 597088
rect 399678 597032 417250 597088
rect 417306 597032 417374 597088
rect 417430 597032 417498 597088
rect 417554 597032 417622 597088
rect 417678 597032 435250 597088
rect 435306 597032 435374 597088
rect 435430 597032 435498 597088
rect 435554 597032 435622 597088
rect 435678 597032 453250 597088
rect 453306 597032 453374 597088
rect 453430 597032 453498 597088
rect 453554 597032 453622 597088
rect 453678 597032 471250 597088
rect 471306 597032 471374 597088
rect 471430 597032 471498 597088
rect 471554 597032 471622 597088
rect 471678 597032 489250 597088
rect 489306 597032 489374 597088
rect 489430 597032 489498 597088
rect 489554 597032 489622 597088
rect 489678 597032 507250 597088
rect 507306 597032 507374 597088
rect 507430 597032 507498 597088
rect 507554 597032 507622 597088
rect 507678 597032 525250 597088
rect 525306 597032 525374 597088
rect 525430 597032 525498 597088
rect 525554 597032 525622 597088
rect 525678 597032 543250 597088
rect 543306 597032 543374 597088
rect 543430 597032 543498 597088
rect 543554 597032 543622 597088
rect 543678 597032 561250 597088
rect 561306 597032 561374 597088
rect 561430 597032 561498 597088
rect 561554 597032 561622 597088
rect 561678 597032 579250 597088
rect 579306 597032 579374 597088
rect 579430 597032 579498 597088
rect 579554 597032 579622 597088
rect 579678 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect -956 596964 597020 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 3250 596964
rect 3306 596908 3374 596964
rect 3430 596908 3498 596964
rect 3554 596908 3622 596964
rect 3678 596908 21250 596964
rect 21306 596908 21374 596964
rect 21430 596908 21498 596964
rect 21554 596908 21622 596964
rect 21678 596908 39250 596964
rect 39306 596908 39374 596964
rect 39430 596908 39498 596964
rect 39554 596908 39622 596964
rect 39678 596908 57250 596964
rect 57306 596908 57374 596964
rect 57430 596908 57498 596964
rect 57554 596908 57622 596964
rect 57678 596908 75250 596964
rect 75306 596908 75374 596964
rect 75430 596908 75498 596964
rect 75554 596908 75622 596964
rect 75678 596908 93250 596964
rect 93306 596908 93374 596964
rect 93430 596908 93498 596964
rect 93554 596908 93622 596964
rect 93678 596908 111250 596964
rect 111306 596908 111374 596964
rect 111430 596908 111498 596964
rect 111554 596908 111622 596964
rect 111678 596908 129250 596964
rect 129306 596908 129374 596964
rect 129430 596908 129498 596964
rect 129554 596908 129622 596964
rect 129678 596908 147250 596964
rect 147306 596908 147374 596964
rect 147430 596908 147498 596964
rect 147554 596908 147622 596964
rect 147678 596908 165250 596964
rect 165306 596908 165374 596964
rect 165430 596908 165498 596964
rect 165554 596908 165622 596964
rect 165678 596908 183250 596964
rect 183306 596908 183374 596964
rect 183430 596908 183498 596964
rect 183554 596908 183622 596964
rect 183678 596908 201250 596964
rect 201306 596908 201374 596964
rect 201430 596908 201498 596964
rect 201554 596908 201622 596964
rect 201678 596908 219250 596964
rect 219306 596908 219374 596964
rect 219430 596908 219498 596964
rect 219554 596908 219622 596964
rect 219678 596908 237250 596964
rect 237306 596908 237374 596964
rect 237430 596908 237498 596964
rect 237554 596908 237622 596964
rect 237678 596908 255250 596964
rect 255306 596908 255374 596964
rect 255430 596908 255498 596964
rect 255554 596908 255622 596964
rect 255678 596908 273250 596964
rect 273306 596908 273374 596964
rect 273430 596908 273498 596964
rect 273554 596908 273622 596964
rect 273678 596908 291250 596964
rect 291306 596908 291374 596964
rect 291430 596908 291498 596964
rect 291554 596908 291622 596964
rect 291678 596908 309250 596964
rect 309306 596908 309374 596964
rect 309430 596908 309498 596964
rect 309554 596908 309622 596964
rect 309678 596908 327250 596964
rect 327306 596908 327374 596964
rect 327430 596908 327498 596964
rect 327554 596908 327622 596964
rect 327678 596908 345250 596964
rect 345306 596908 345374 596964
rect 345430 596908 345498 596964
rect 345554 596908 345622 596964
rect 345678 596908 363250 596964
rect 363306 596908 363374 596964
rect 363430 596908 363498 596964
rect 363554 596908 363622 596964
rect 363678 596908 381250 596964
rect 381306 596908 381374 596964
rect 381430 596908 381498 596964
rect 381554 596908 381622 596964
rect 381678 596908 399250 596964
rect 399306 596908 399374 596964
rect 399430 596908 399498 596964
rect 399554 596908 399622 596964
rect 399678 596908 417250 596964
rect 417306 596908 417374 596964
rect 417430 596908 417498 596964
rect 417554 596908 417622 596964
rect 417678 596908 435250 596964
rect 435306 596908 435374 596964
rect 435430 596908 435498 596964
rect 435554 596908 435622 596964
rect 435678 596908 453250 596964
rect 453306 596908 453374 596964
rect 453430 596908 453498 596964
rect 453554 596908 453622 596964
rect 453678 596908 471250 596964
rect 471306 596908 471374 596964
rect 471430 596908 471498 596964
rect 471554 596908 471622 596964
rect 471678 596908 489250 596964
rect 489306 596908 489374 596964
rect 489430 596908 489498 596964
rect 489554 596908 489622 596964
rect 489678 596908 507250 596964
rect 507306 596908 507374 596964
rect 507430 596908 507498 596964
rect 507554 596908 507622 596964
rect 507678 596908 525250 596964
rect 525306 596908 525374 596964
rect 525430 596908 525498 596964
rect 525554 596908 525622 596964
rect 525678 596908 543250 596964
rect 543306 596908 543374 596964
rect 543430 596908 543498 596964
rect 543554 596908 543622 596964
rect 543678 596908 561250 596964
rect 561306 596908 561374 596964
rect 561430 596908 561498 596964
rect 561554 596908 561622 596964
rect 561678 596908 579250 596964
rect 579306 596908 579374 596964
rect 579430 596908 579498 596964
rect 579554 596908 579622 596964
rect 579678 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect -956 596840 597020 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 3250 596840
rect 3306 596784 3374 596840
rect 3430 596784 3498 596840
rect 3554 596784 3622 596840
rect 3678 596784 21250 596840
rect 21306 596784 21374 596840
rect 21430 596784 21498 596840
rect 21554 596784 21622 596840
rect 21678 596784 39250 596840
rect 39306 596784 39374 596840
rect 39430 596784 39498 596840
rect 39554 596784 39622 596840
rect 39678 596784 57250 596840
rect 57306 596784 57374 596840
rect 57430 596784 57498 596840
rect 57554 596784 57622 596840
rect 57678 596784 75250 596840
rect 75306 596784 75374 596840
rect 75430 596784 75498 596840
rect 75554 596784 75622 596840
rect 75678 596784 93250 596840
rect 93306 596784 93374 596840
rect 93430 596784 93498 596840
rect 93554 596784 93622 596840
rect 93678 596784 111250 596840
rect 111306 596784 111374 596840
rect 111430 596784 111498 596840
rect 111554 596784 111622 596840
rect 111678 596784 129250 596840
rect 129306 596784 129374 596840
rect 129430 596784 129498 596840
rect 129554 596784 129622 596840
rect 129678 596784 147250 596840
rect 147306 596784 147374 596840
rect 147430 596784 147498 596840
rect 147554 596784 147622 596840
rect 147678 596784 165250 596840
rect 165306 596784 165374 596840
rect 165430 596784 165498 596840
rect 165554 596784 165622 596840
rect 165678 596784 183250 596840
rect 183306 596784 183374 596840
rect 183430 596784 183498 596840
rect 183554 596784 183622 596840
rect 183678 596784 201250 596840
rect 201306 596784 201374 596840
rect 201430 596784 201498 596840
rect 201554 596784 201622 596840
rect 201678 596784 219250 596840
rect 219306 596784 219374 596840
rect 219430 596784 219498 596840
rect 219554 596784 219622 596840
rect 219678 596784 237250 596840
rect 237306 596784 237374 596840
rect 237430 596784 237498 596840
rect 237554 596784 237622 596840
rect 237678 596784 255250 596840
rect 255306 596784 255374 596840
rect 255430 596784 255498 596840
rect 255554 596784 255622 596840
rect 255678 596784 273250 596840
rect 273306 596784 273374 596840
rect 273430 596784 273498 596840
rect 273554 596784 273622 596840
rect 273678 596784 291250 596840
rect 291306 596784 291374 596840
rect 291430 596784 291498 596840
rect 291554 596784 291622 596840
rect 291678 596784 309250 596840
rect 309306 596784 309374 596840
rect 309430 596784 309498 596840
rect 309554 596784 309622 596840
rect 309678 596784 327250 596840
rect 327306 596784 327374 596840
rect 327430 596784 327498 596840
rect 327554 596784 327622 596840
rect 327678 596784 345250 596840
rect 345306 596784 345374 596840
rect 345430 596784 345498 596840
rect 345554 596784 345622 596840
rect 345678 596784 363250 596840
rect 363306 596784 363374 596840
rect 363430 596784 363498 596840
rect 363554 596784 363622 596840
rect 363678 596784 381250 596840
rect 381306 596784 381374 596840
rect 381430 596784 381498 596840
rect 381554 596784 381622 596840
rect 381678 596784 399250 596840
rect 399306 596784 399374 596840
rect 399430 596784 399498 596840
rect 399554 596784 399622 596840
rect 399678 596784 417250 596840
rect 417306 596784 417374 596840
rect 417430 596784 417498 596840
rect 417554 596784 417622 596840
rect 417678 596784 435250 596840
rect 435306 596784 435374 596840
rect 435430 596784 435498 596840
rect 435554 596784 435622 596840
rect 435678 596784 453250 596840
rect 453306 596784 453374 596840
rect 453430 596784 453498 596840
rect 453554 596784 453622 596840
rect 453678 596784 471250 596840
rect 471306 596784 471374 596840
rect 471430 596784 471498 596840
rect 471554 596784 471622 596840
rect 471678 596784 489250 596840
rect 489306 596784 489374 596840
rect 489430 596784 489498 596840
rect 489554 596784 489622 596840
rect 489678 596784 507250 596840
rect 507306 596784 507374 596840
rect 507430 596784 507498 596840
rect 507554 596784 507622 596840
rect 507678 596784 525250 596840
rect 525306 596784 525374 596840
rect 525430 596784 525498 596840
rect 525554 596784 525622 596840
rect 525678 596784 543250 596840
rect 543306 596784 543374 596840
rect 543430 596784 543498 596840
rect 543554 596784 543622 596840
rect 543678 596784 561250 596840
rect 561306 596784 561374 596840
rect 561430 596784 561498 596840
rect 561554 596784 561622 596840
rect 561678 596784 579250 596840
rect 579306 596784 579374 596840
rect 579430 596784 579498 596840
rect 579554 596784 579622 596840
rect 579678 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect -956 596688 597020 596784
rect -1916 586350 597980 586446
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 6970 586350
rect 7026 586294 7094 586350
rect 7150 586294 7218 586350
rect 7274 586294 7342 586350
rect 7398 586294 24970 586350
rect 25026 586294 25094 586350
rect 25150 586294 25218 586350
rect 25274 586294 25342 586350
rect 25398 586294 42970 586350
rect 43026 586294 43094 586350
rect 43150 586294 43218 586350
rect 43274 586294 43342 586350
rect 43398 586294 60970 586350
rect 61026 586294 61094 586350
rect 61150 586294 61218 586350
rect 61274 586294 61342 586350
rect 61398 586294 78970 586350
rect 79026 586294 79094 586350
rect 79150 586294 79218 586350
rect 79274 586294 79342 586350
rect 79398 586294 96970 586350
rect 97026 586294 97094 586350
rect 97150 586294 97218 586350
rect 97274 586294 97342 586350
rect 97398 586294 114970 586350
rect 115026 586294 115094 586350
rect 115150 586294 115218 586350
rect 115274 586294 115342 586350
rect 115398 586294 132970 586350
rect 133026 586294 133094 586350
rect 133150 586294 133218 586350
rect 133274 586294 133342 586350
rect 133398 586294 150970 586350
rect 151026 586294 151094 586350
rect 151150 586294 151218 586350
rect 151274 586294 151342 586350
rect 151398 586294 168970 586350
rect 169026 586294 169094 586350
rect 169150 586294 169218 586350
rect 169274 586294 169342 586350
rect 169398 586294 186970 586350
rect 187026 586294 187094 586350
rect 187150 586294 187218 586350
rect 187274 586294 187342 586350
rect 187398 586294 204970 586350
rect 205026 586294 205094 586350
rect 205150 586294 205218 586350
rect 205274 586294 205342 586350
rect 205398 586294 222970 586350
rect 223026 586294 223094 586350
rect 223150 586294 223218 586350
rect 223274 586294 223342 586350
rect 223398 586294 240970 586350
rect 241026 586294 241094 586350
rect 241150 586294 241218 586350
rect 241274 586294 241342 586350
rect 241398 586294 258970 586350
rect 259026 586294 259094 586350
rect 259150 586294 259218 586350
rect 259274 586294 259342 586350
rect 259398 586294 276970 586350
rect 277026 586294 277094 586350
rect 277150 586294 277218 586350
rect 277274 586294 277342 586350
rect 277398 586294 294970 586350
rect 295026 586294 295094 586350
rect 295150 586294 295218 586350
rect 295274 586294 295342 586350
rect 295398 586294 312970 586350
rect 313026 586294 313094 586350
rect 313150 586294 313218 586350
rect 313274 586294 313342 586350
rect 313398 586294 330970 586350
rect 331026 586294 331094 586350
rect 331150 586294 331218 586350
rect 331274 586294 331342 586350
rect 331398 586294 348970 586350
rect 349026 586294 349094 586350
rect 349150 586294 349218 586350
rect 349274 586294 349342 586350
rect 349398 586294 366970 586350
rect 367026 586294 367094 586350
rect 367150 586294 367218 586350
rect 367274 586294 367342 586350
rect 367398 586294 384970 586350
rect 385026 586294 385094 586350
rect 385150 586294 385218 586350
rect 385274 586294 385342 586350
rect 385398 586294 402970 586350
rect 403026 586294 403094 586350
rect 403150 586294 403218 586350
rect 403274 586294 403342 586350
rect 403398 586294 420970 586350
rect 421026 586294 421094 586350
rect 421150 586294 421218 586350
rect 421274 586294 421342 586350
rect 421398 586294 438970 586350
rect 439026 586294 439094 586350
rect 439150 586294 439218 586350
rect 439274 586294 439342 586350
rect 439398 586294 456970 586350
rect 457026 586294 457094 586350
rect 457150 586294 457218 586350
rect 457274 586294 457342 586350
rect 457398 586294 474970 586350
rect 475026 586294 475094 586350
rect 475150 586294 475218 586350
rect 475274 586294 475342 586350
rect 475398 586294 492970 586350
rect 493026 586294 493094 586350
rect 493150 586294 493218 586350
rect 493274 586294 493342 586350
rect 493398 586294 510970 586350
rect 511026 586294 511094 586350
rect 511150 586294 511218 586350
rect 511274 586294 511342 586350
rect 511398 586294 528970 586350
rect 529026 586294 529094 586350
rect 529150 586294 529218 586350
rect 529274 586294 529342 586350
rect 529398 586294 546970 586350
rect 547026 586294 547094 586350
rect 547150 586294 547218 586350
rect 547274 586294 547342 586350
rect 547398 586294 564970 586350
rect 565026 586294 565094 586350
rect 565150 586294 565218 586350
rect 565274 586294 565342 586350
rect 565398 586294 582970 586350
rect 583026 586294 583094 586350
rect 583150 586294 583218 586350
rect 583274 586294 583342 586350
rect 583398 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect -1916 586226 597980 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 6970 586226
rect 7026 586170 7094 586226
rect 7150 586170 7218 586226
rect 7274 586170 7342 586226
rect 7398 586170 24970 586226
rect 25026 586170 25094 586226
rect 25150 586170 25218 586226
rect 25274 586170 25342 586226
rect 25398 586170 42970 586226
rect 43026 586170 43094 586226
rect 43150 586170 43218 586226
rect 43274 586170 43342 586226
rect 43398 586170 60970 586226
rect 61026 586170 61094 586226
rect 61150 586170 61218 586226
rect 61274 586170 61342 586226
rect 61398 586170 78970 586226
rect 79026 586170 79094 586226
rect 79150 586170 79218 586226
rect 79274 586170 79342 586226
rect 79398 586170 96970 586226
rect 97026 586170 97094 586226
rect 97150 586170 97218 586226
rect 97274 586170 97342 586226
rect 97398 586170 114970 586226
rect 115026 586170 115094 586226
rect 115150 586170 115218 586226
rect 115274 586170 115342 586226
rect 115398 586170 132970 586226
rect 133026 586170 133094 586226
rect 133150 586170 133218 586226
rect 133274 586170 133342 586226
rect 133398 586170 150970 586226
rect 151026 586170 151094 586226
rect 151150 586170 151218 586226
rect 151274 586170 151342 586226
rect 151398 586170 168970 586226
rect 169026 586170 169094 586226
rect 169150 586170 169218 586226
rect 169274 586170 169342 586226
rect 169398 586170 186970 586226
rect 187026 586170 187094 586226
rect 187150 586170 187218 586226
rect 187274 586170 187342 586226
rect 187398 586170 204970 586226
rect 205026 586170 205094 586226
rect 205150 586170 205218 586226
rect 205274 586170 205342 586226
rect 205398 586170 222970 586226
rect 223026 586170 223094 586226
rect 223150 586170 223218 586226
rect 223274 586170 223342 586226
rect 223398 586170 240970 586226
rect 241026 586170 241094 586226
rect 241150 586170 241218 586226
rect 241274 586170 241342 586226
rect 241398 586170 258970 586226
rect 259026 586170 259094 586226
rect 259150 586170 259218 586226
rect 259274 586170 259342 586226
rect 259398 586170 276970 586226
rect 277026 586170 277094 586226
rect 277150 586170 277218 586226
rect 277274 586170 277342 586226
rect 277398 586170 294970 586226
rect 295026 586170 295094 586226
rect 295150 586170 295218 586226
rect 295274 586170 295342 586226
rect 295398 586170 312970 586226
rect 313026 586170 313094 586226
rect 313150 586170 313218 586226
rect 313274 586170 313342 586226
rect 313398 586170 330970 586226
rect 331026 586170 331094 586226
rect 331150 586170 331218 586226
rect 331274 586170 331342 586226
rect 331398 586170 348970 586226
rect 349026 586170 349094 586226
rect 349150 586170 349218 586226
rect 349274 586170 349342 586226
rect 349398 586170 366970 586226
rect 367026 586170 367094 586226
rect 367150 586170 367218 586226
rect 367274 586170 367342 586226
rect 367398 586170 384970 586226
rect 385026 586170 385094 586226
rect 385150 586170 385218 586226
rect 385274 586170 385342 586226
rect 385398 586170 402970 586226
rect 403026 586170 403094 586226
rect 403150 586170 403218 586226
rect 403274 586170 403342 586226
rect 403398 586170 420970 586226
rect 421026 586170 421094 586226
rect 421150 586170 421218 586226
rect 421274 586170 421342 586226
rect 421398 586170 438970 586226
rect 439026 586170 439094 586226
rect 439150 586170 439218 586226
rect 439274 586170 439342 586226
rect 439398 586170 456970 586226
rect 457026 586170 457094 586226
rect 457150 586170 457218 586226
rect 457274 586170 457342 586226
rect 457398 586170 474970 586226
rect 475026 586170 475094 586226
rect 475150 586170 475218 586226
rect 475274 586170 475342 586226
rect 475398 586170 492970 586226
rect 493026 586170 493094 586226
rect 493150 586170 493218 586226
rect 493274 586170 493342 586226
rect 493398 586170 510970 586226
rect 511026 586170 511094 586226
rect 511150 586170 511218 586226
rect 511274 586170 511342 586226
rect 511398 586170 528970 586226
rect 529026 586170 529094 586226
rect 529150 586170 529218 586226
rect 529274 586170 529342 586226
rect 529398 586170 546970 586226
rect 547026 586170 547094 586226
rect 547150 586170 547218 586226
rect 547274 586170 547342 586226
rect 547398 586170 564970 586226
rect 565026 586170 565094 586226
rect 565150 586170 565218 586226
rect 565274 586170 565342 586226
rect 565398 586170 582970 586226
rect 583026 586170 583094 586226
rect 583150 586170 583218 586226
rect 583274 586170 583342 586226
rect 583398 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect -1916 586102 597980 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 6970 586102
rect 7026 586046 7094 586102
rect 7150 586046 7218 586102
rect 7274 586046 7342 586102
rect 7398 586046 24970 586102
rect 25026 586046 25094 586102
rect 25150 586046 25218 586102
rect 25274 586046 25342 586102
rect 25398 586046 42970 586102
rect 43026 586046 43094 586102
rect 43150 586046 43218 586102
rect 43274 586046 43342 586102
rect 43398 586046 60970 586102
rect 61026 586046 61094 586102
rect 61150 586046 61218 586102
rect 61274 586046 61342 586102
rect 61398 586046 78970 586102
rect 79026 586046 79094 586102
rect 79150 586046 79218 586102
rect 79274 586046 79342 586102
rect 79398 586046 96970 586102
rect 97026 586046 97094 586102
rect 97150 586046 97218 586102
rect 97274 586046 97342 586102
rect 97398 586046 114970 586102
rect 115026 586046 115094 586102
rect 115150 586046 115218 586102
rect 115274 586046 115342 586102
rect 115398 586046 132970 586102
rect 133026 586046 133094 586102
rect 133150 586046 133218 586102
rect 133274 586046 133342 586102
rect 133398 586046 150970 586102
rect 151026 586046 151094 586102
rect 151150 586046 151218 586102
rect 151274 586046 151342 586102
rect 151398 586046 168970 586102
rect 169026 586046 169094 586102
rect 169150 586046 169218 586102
rect 169274 586046 169342 586102
rect 169398 586046 186970 586102
rect 187026 586046 187094 586102
rect 187150 586046 187218 586102
rect 187274 586046 187342 586102
rect 187398 586046 204970 586102
rect 205026 586046 205094 586102
rect 205150 586046 205218 586102
rect 205274 586046 205342 586102
rect 205398 586046 222970 586102
rect 223026 586046 223094 586102
rect 223150 586046 223218 586102
rect 223274 586046 223342 586102
rect 223398 586046 240970 586102
rect 241026 586046 241094 586102
rect 241150 586046 241218 586102
rect 241274 586046 241342 586102
rect 241398 586046 258970 586102
rect 259026 586046 259094 586102
rect 259150 586046 259218 586102
rect 259274 586046 259342 586102
rect 259398 586046 276970 586102
rect 277026 586046 277094 586102
rect 277150 586046 277218 586102
rect 277274 586046 277342 586102
rect 277398 586046 294970 586102
rect 295026 586046 295094 586102
rect 295150 586046 295218 586102
rect 295274 586046 295342 586102
rect 295398 586046 312970 586102
rect 313026 586046 313094 586102
rect 313150 586046 313218 586102
rect 313274 586046 313342 586102
rect 313398 586046 330970 586102
rect 331026 586046 331094 586102
rect 331150 586046 331218 586102
rect 331274 586046 331342 586102
rect 331398 586046 348970 586102
rect 349026 586046 349094 586102
rect 349150 586046 349218 586102
rect 349274 586046 349342 586102
rect 349398 586046 366970 586102
rect 367026 586046 367094 586102
rect 367150 586046 367218 586102
rect 367274 586046 367342 586102
rect 367398 586046 384970 586102
rect 385026 586046 385094 586102
rect 385150 586046 385218 586102
rect 385274 586046 385342 586102
rect 385398 586046 402970 586102
rect 403026 586046 403094 586102
rect 403150 586046 403218 586102
rect 403274 586046 403342 586102
rect 403398 586046 420970 586102
rect 421026 586046 421094 586102
rect 421150 586046 421218 586102
rect 421274 586046 421342 586102
rect 421398 586046 438970 586102
rect 439026 586046 439094 586102
rect 439150 586046 439218 586102
rect 439274 586046 439342 586102
rect 439398 586046 456970 586102
rect 457026 586046 457094 586102
rect 457150 586046 457218 586102
rect 457274 586046 457342 586102
rect 457398 586046 474970 586102
rect 475026 586046 475094 586102
rect 475150 586046 475218 586102
rect 475274 586046 475342 586102
rect 475398 586046 492970 586102
rect 493026 586046 493094 586102
rect 493150 586046 493218 586102
rect 493274 586046 493342 586102
rect 493398 586046 510970 586102
rect 511026 586046 511094 586102
rect 511150 586046 511218 586102
rect 511274 586046 511342 586102
rect 511398 586046 528970 586102
rect 529026 586046 529094 586102
rect 529150 586046 529218 586102
rect 529274 586046 529342 586102
rect 529398 586046 546970 586102
rect 547026 586046 547094 586102
rect 547150 586046 547218 586102
rect 547274 586046 547342 586102
rect 547398 586046 564970 586102
rect 565026 586046 565094 586102
rect 565150 586046 565218 586102
rect 565274 586046 565342 586102
rect 565398 586046 582970 586102
rect 583026 586046 583094 586102
rect 583150 586046 583218 586102
rect 583274 586046 583342 586102
rect 583398 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect -1916 585978 597980 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 6970 585978
rect 7026 585922 7094 585978
rect 7150 585922 7218 585978
rect 7274 585922 7342 585978
rect 7398 585922 24970 585978
rect 25026 585922 25094 585978
rect 25150 585922 25218 585978
rect 25274 585922 25342 585978
rect 25398 585922 42970 585978
rect 43026 585922 43094 585978
rect 43150 585922 43218 585978
rect 43274 585922 43342 585978
rect 43398 585922 60970 585978
rect 61026 585922 61094 585978
rect 61150 585922 61218 585978
rect 61274 585922 61342 585978
rect 61398 585922 78970 585978
rect 79026 585922 79094 585978
rect 79150 585922 79218 585978
rect 79274 585922 79342 585978
rect 79398 585922 96970 585978
rect 97026 585922 97094 585978
rect 97150 585922 97218 585978
rect 97274 585922 97342 585978
rect 97398 585922 114970 585978
rect 115026 585922 115094 585978
rect 115150 585922 115218 585978
rect 115274 585922 115342 585978
rect 115398 585922 132970 585978
rect 133026 585922 133094 585978
rect 133150 585922 133218 585978
rect 133274 585922 133342 585978
rect 133398 585922 150970 585978
rect 151026 585922 151094 585978
rect 151150 585922 151218 585978
rect 151274 585922 151342 585978
rect 151398 585922 168970 585978
rect 169026 585922 169094 585978
rect 169150 585922 169218 585978
rect 169274 585922 169342 585978
rect 169398 585922 186970 585978
rect 187026 585922 187094 585978
rect 187150 585922 187218 585978
rect 187274 585922 187342 585978
rect 187398 585922 204970 585978
rect 205026 585922 205094 585978
rect 205150 585922 205218 585978
rect 205274 585922 205342 585978
rect 205398 585922 222970 585978
rect 223026 585922 223094 585978
rect 223150 585922 223218 585978
rect 223274 585922 223342 585978
rect 223398 585922 240970 585978
rect 241026 585922 241094 585978
rect 241150 585922 241218 585978
rect 241274 585922 241342 585978
rect 241398 585922 258970 585978
rect 259026 585922 259094 585978
rect 259150 585922 259218 585978
rect 259274 585922 259342 585978
rect 259398 585922 276970 585978
rect 277026 585922 277094 585978
rect 277150 585922 277218 585978
rect 277274 585922 277342 585978
rect 277398 585922 294970 585978
rect 295026 585922 295094 585978
rect 295150 585922 295218 585978
rect 295274 585922 295342 585978
rect 295398 585922 312970 585978
rect 313026 585922 313094 585978
rect 313150 585922 313218 585978
rect 313274 585922 313342 585978
rect 313398 585922 330970 585978
rect 331026 585922 331094 585978
rect 331150 585922 331218 585978
rect 331274 585922 331342 585978
rect 331398 585922 348970 585978
rect 349026 585922 349094 585978
rect 349150 585922 349218 585978
rect 349274 585922 349342 585978
rect 349398 585922 366970 585978
rect 367026 585922 367094 585978
rect 367150 585922 367218 585978
rect 367274 585922 367342 585978
rect 367398 585922 384970 585978
rect 385026 585922 385094 585978
rect 385150 585922 385218 585978
rect 385274 585922 385342 585978
rect 385398 585922 402970 585978
rect 403026 585922 403094 585978
rect 403150 585922 403218 585978
rect 403274 585922 403342 585978
rect 403398 585922 420970 585978
rect 421026 585922 421094 585978
rect 421150 585922 421218 585978
rect 421274 585922 421342 585978
rect 421398 585922 438970 585978
rect 439026 585922 439094 585978
rect 439150 585922 439218 585978
rect 439274 585922 439342 585978
rect 439398 585922 456970 585978
rect 457026 585922 457094 585978
rect 457150 585922 457218 585978
rect 457274 585922 457342 585978
rect 457398 585922 474970 585978
rect 475026 585922 475094 585978
rect 475150 585922 475218 585978
rect 475274 585922 475342 585978
rect 475398 585922 492970 585978
rect 493026 585922 493094 585978
rect 493150 585922 493218 585978
rect 493274 585922 493342 585978
rect 493398 585922 510970 585978
rect 511026 585922 511094 585978
rect 511150 585922 511218 585978
rect 511274 585922 511342 585978
rect 511398 585922 528970 585978
rect 529026 585922 529094 585978
rect 529150 585922 529218 585978
rect 529274 585922 529342 585978
rect 529398 585922 546970 585978
rect 547026 585922 547094 585978
rect 547150 585922 547218 585978
rect 547274 585922 547342 585978
rect 547398 585922 564970 585978
rect 565026 585922 565094 585978
rect 565150 585922 565218 585978
rect 565274 585922 565342 585978
rect 565398 585922 582970 585978
rect 583026 585922 583094 585978
rect 583150 585922 583218 585978
rect 583274 585922 583342 585978
rect 583398 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect -1916 585826 597980 585922
rect -1916 580350 597980 580446
rect -1916 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 3250 580350
rect 3306 580294 3374 580350
rect 3430 580294 3498 580350
rect 3554 580294 3622 580350
rect 3678 580294 21250 580350
rect 21306 580294 21374 580350
rect 21430 580294 21498 580350
rect 21554 580294 21622 580350
rect 21678 580294 39250 580350
rect 39306 580294 39374 580350
rect 39430 580294 39498 580350
rect 39554 580294 39622 580350
rect 39678 580294 57250 580350
rect 57306 580294 57374 580350
rect 57430 580294 57498 580350
rect 57554 580294 57622 580350
rect 57678 580294 75250 580350
rect 75306 580294 75374 580350
rect 75430 580294 75498 580350
rect 75554 580294 75622 580350
rect 75678 580294 93250 580350
rect 93306 580294 93374 580350
rect 93430 580294 93498 580350
rect 93554 580294 93622 580350
rect 93678 580294 111250 580350
rect 111306 580294 111374 580350
rect 111430 580294 111498 580350
rect 111554 580294 111622 580350
rect 111678 580294 129250 580350
rect 129306 580294 129374 580350
rect 129430 580294 129498 580350
rect 129554 580294 129622 580350
rect 129678 580294 147250 580350
rect 147306 580294 147374 580350
rect 147430 580294 147498 580350
rect 147554 580294 147622 580350
rect 147678 580294 165250 580350
rect 165306 580294 165374 580350
rect 165430 580294 165498 580350
rect 165554 580294 165622 580350
rect 165678 580294 183250 580350
rect 183306 580294 183374 580350
rect 183430 580294 183498 580350
rect 183554 580294 183622 580350
rect 183678 580294 201250 580350
rect 201306 580294 201374 580350
rect 201430 580294 201498 580350
rect 201554 580294 201622 580350
rect 201678 580294 219250 580350
rect 219306 580294 219374 580350
rect 219430 580294 219498 580350
rect 219554 580294 219622 580350
rect 219678 580294 237250 580350
rect 237306 580294 237374 580350
rect 237430 580294 237498 580350
rect 237554 580294 237622 580350
rect 237678 580294 255250 580350
rect 255306 580294 255374 580350
rect 255430 580294 255498 580350
rect 255554 580294 255622 580350
rect 255678 580294 273250 580350
rect 273306 580294 273374 580350
rect 273430 580294 273498 580350
rect 273554 580294 273622 580350
rect 273678 580294 291250 580350
rect 291306 580294 291374 580350
rect 291430 580294 291498 580350
rect 291554 580294 291622 580350
rect 291678 580294 309250 580350
rect 309306 580294 309374 580350
rect 309430 580294 309498 580350
rect 309554 580294 309622 580350
rect 309678 580294 327250 580350
rect 327306 580294 327374 580350
rect 327430 580294 327498 580350
rect 327554 580294 327622 580350
rect 327678 580294 345250 580350
rect 345306 580294 345374 580350
rect 345430 580294 345498 580350
rect 345554 580294 345622 580350
rect 345678 580294 363250 580350
rect 363306 580294 363374 580350
rect 363430 580294 363498 580350
rect 363554 580294 363622 580350
rect 363678 580294 381250 580350
rect 381306 580294 381374 580350
rect 381430 580294 381498 580350
rect 381554 580294 381622 580350
rect 381678 580294 399250 580350
rect 399306 580294 399374 580350
rect 399430 580294 399498 580350
rect 399554 580294 399622 580350
rect 399678 580294 417250 580350
rect 417306 580294 417374 580350
rect 417430 580294 417498 580350
rect 417554 580294 417622 580350
rect 417678 580294 435250 580350
rect 435306 580294 435374 580350
rect 435430 580294 435498 580350
rect 435554 580294 435622 580350
rect 435678 580294 453250 580350
rect 453306 580294 453374 580350
rect 453430 580294 453498 580350
rect 453554 580294 453622 580350
rect 453678 580294 471250 580350
rect 471306 580294 471374 580350
rect 471430 580294 471498 580350
rect 471554 580294 471622 580350
rect 471678 580294 489250 580350
rect 489306 580294 489374 580350
rect 489430 580294 489498 580350
rect 489554 580294 489622 580350
rect 489678 580294 507250 580350
rect 507306 580294 507374 580350
rect 507430 580294 507498 580350
rect 507554 580294 507622 580350
rect 507678 580294 525250 580350
rect 525306 580294 525374 580350
rect 525430 580294 525498 580350
rect 525554 580294 525622 580350
rect 525678 580294 543250 580350
rect 543306 580294 543374 580350
rect 543430 580294 543498 580350
rect 543554 580294 543622 580350
rect 543678 580294 561250 580350
rect 561306 580294 561374 580350
rect 561430 580294 561498 580350
rect 561554 580294 561622 580350
rect 561678 580294 579250 580350
rect 579306 580294 579374 580350
rect 579430 580294 579498 580350
rect 579554 580294 579622 580350
rect 579678 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597980 580350
rect -1916 580226 597980 580294
rect -1916 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 3250 580226
rect 3306 580170 3374 580226
rect 3430 580170 3498 580226
rect 3554 580170 3622 580226
rect 3678 580170 21250 580226
rect 21306 580170 21374 580226
rect 21430 580170 21498 580226
rect 21554 580170 21622 580226
rect 21678 580170 39250 580226
rect 39306 580170 39374 580226
rect 39430 580170 39498 580226
rect 39554 580170 39622 580226
rect 39678 580170 57250 580226
rect 57306 580170 57374 580226
rect 57430 580170 57498 580226
rect 57554 580170 57622 580226
rect 57678 580170 75250 580226
rect 75306 580170 75374 580226
rect 75430 580170 75498 580226
rect 75554 580170 75622 580226
rect 75678 580170 93250 580226
rect 93306 580170 93374 580226
rect 93430 580170 93498 580226
rect 93554 580170 93622 580226
rect 93678 580170 111250 580226
rect 111306 580170 111374 580226
rect 111430 580170 111498 580226
rect 111554 580170 111622 580226
rect 111678 580170 129250 580226
rect 129306 580170 129374 580226
rect 129430 580170 129498 580226
rect 129554 580170 129622 580226
rect 129678 580170 147250 580226
rect 147306 580170 147374 580226
rect 147430 580170 147498 580226
rect 147554 580170 147622 580226
rect 147678 580170 165250 580226
rect 165306 580170 165374 580226
rect 165430 580170 165498 580226
rect 165554 580170 165622 580226
rect 165678 580170 183250 580226
rect 183306 580170 183374 580226
rect 183430 580170 183498 580226
rect 183554 580170 183622 580226
rect 183678 580170 201250 580226
rect 201306 580170 201374 580226
rect 201430 580170 201498 580226
rect 201554 580170 201622 580226
rect 201678 580170 219250 580226
rect 219306 580170 219374 580226
rect 219430 580170 219498 580226
rect 219554 580170 219622 580226
rect 219678 580170 237250 580226
rect 237306 580170 237374 580226
rect 237430 580170 237498 580226
rect 237554 580170 237622 580226
rect 237678 580170 255250 580226
rect 255306 580170 255374 580226
rect 255430 580170 255498 580226
rect 255554 580170 255622 580226
rect 255678 580170 273250 580226
rect 273306 580170 273374 580226
rect 273430 580170 273498 580226
rect 273554 580170 273622 580226
rect 273678 580170 291250 580226
rect 291306 580170 291374 580226
rect 291430 580170 291498 580226
rect 291554 580170 291622 580226
rect 291678 580170 309250 580226
rect 309306 580170 309374 580226
rect 309430 580170 309498 580226
rect 309554 580170 309622 580226
rect 309678 580170 327250 580226
rect 327306 580170 327374 580226
rect 327430 580170 327498 580226
rect 327554 580170 327622 580226
rect 327678 580170 345250 580226
rect 345306 580170 345374 580226
rect 345430 580170 345498 580226
rect 345554 580170 345622 580226
rect 345678 580170 363250 580226
rect 363306 580170 363374 580226
rect 363430 580170 363498 580226
rect 363554 580170 363622 580226
rect 363678 580170 381250 580226
rect 381306 580170 381374 580226
rect 381430 580170 381498 580226
rect 381554 580170 381622 580226
rect 381678 580170 399250 580226
rect 399306 580170 399374 580226
rect 399430 580170 399498 580226
rect 399554 580170 399622 580226
rect 399678 580170 417250 580226
rect 417306 580170 417374 580226
rect 417430 580170 417498 580226
rect 417554 580170 417622 580226
rect 417678 580170 435250 580226
rect 435306 580170 435374 580226
rect 435430 580170 435498 580226
rect 435554 580170 435622 580226
rect 435678 580170 453250 580226
rect 453306 580170 453374 580226
rect 453430 580170 453498 580226
rect 453554 580170 453622 580226
rect 453678 580170 471250 580226
rect 471306 580170 471374 580226
rect 471430 580170 471498 580226
rect 471554 580170 471622 580226
rect 471678 580170 489250 580226
rect 489306 580170 489374 580226
rect 489430 580170 489498 580226
rect 489554 580170 489622 580226
rect 489678 580170 507250 580226
rect 507306 580170 507374 580226
rect 507430 580170 507498 580226
rect 507554 580170 507622 580226
rect 507678 580170 525250 580226
rect 525306 580170 525374 580226
rect 525430 580170 525498 580226
rect 525554 580170 525622 580226
rect 525678 580170 543250 580226
rect 543306 580170 543374 580226
rect 543430 580170 543498 580226
rect 543554 580170 543622 580226
rect 543678 580170 561250 580226
rect 561306 580170 561374 580226
rect 561430 580170 561498 580226
rect 561554 580170 561622 580226
rect 561678 580170 579250 580226
rect 579306 580170 579374 580226
rect 579430 580170 579498 580226
rect 579554 580170 579622 580226
rect 579678 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597980 580226
rect -1916 580102 597980 580170
rect -1916 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 3250 580102
rect 3306 580046 3374 580102
rect 3430 580046 3498 580102
rect 3554 580046 3622 580102
rect 3678 580046 21250 580102
rect 21306 580046 21374 580102
rect 21430 580046 21498 580102
rect 21554 580046 21622 580102
rect 21678 580046 39250 580102
rect 39306 580046 39374 580102
rect 39430 580046 39498 580102
rect 39554 580046 39622 580102
rect 39678 580046 57250 580102
rect 57306 580046 57374 580102
rect 57430 580046 57498 580102
rect 57554 580046 57622 580102
rect 57678 580046 75250 580102
rect 75306 580046 75374 580102
rect 75430 580046 75498 580102
rect 75554 580046 75622 580102
rect 75678 580046 93250 580102
rect 93306 580046 93374 580102
rect 93430 580046 93498 580102
rect 93554 580046 93622 580102
rect 93678 580046 111250 580102
rect 111306 580046 111374 580102
rect 111430 580046 111498 580102
rect 111554 580046 111622 580102
rect 111678 580046 129250 580102
rect 129306 580046 129374 580102
rect 129430 580046 129498 580102
rect 129554 580046 129622 580102
rect 129678 580046 147250 580102
rect 147306 580046 147374 580102
rect 147430 580046 147498 580102
rect 147554 580046 147622 580102
rect 147678 580046 165250 580102
rect 165306 580046 165374 580102
rect 165430 580046 165498 580102
rect 165554 580046 165622 580102
rect 165678 580046 183250 580102
rect 183306 580046 183374 580102
rect 183430 580046 183498 580102
rect 183554 580046 183622 580102
rect 183678 580046 201250 580102
rect 201306 580046 201374 580102
rect 201430 580046 201498 580102
rect 201554 580046 201622 580102
rect 201678 580046 219250 580102
rect 219306 580046 219374 580102
rect 219430 580046 219498 580102
rect 219554 580046 219622 580102
rect 219678 580046 237250 580102
rect 237306 580046 237374 580102
rect 237430 580046 237498 580102
rect 237554 580046 237622 580102
rect 237678 580046 255250 580102
rect 255306 580046 255374 580102
rect 255430 580046 255498 580102
rect 255554 580046 255622 580102
rect 255678 580046 273250 580102
rect 273306 580046 273374 580102
rect 273430 580046 273498 580102
rect 273554 580046 273622 580102
rect 273678 580046 291250 580102
rect 291306 580046 291374 580102
rect 291430 580046 291498 580102
rect 291554 580046 291622 580102
rect 291678 580046 309250 580102
rect 309306 580046 309374 580102
rect 309430 580046 309498 580102
rect 309554 580046 309622 580102
rect 309678 580046 327250 580102
rect 327306 580046 327374 580102
rect 327430 580046 327498 580102
rect 327554 580046 327622 580102
rect 327678 580046 345250 580102
rect 345306 580046 345374 580102
rect 345430 580046 345498 580102
rect 345554 580046 345622 580102
rect 345678 580046 363250 580102
rect 363306 580046 363374 580102
rect 363430 580046 363498 580102
rect 363554 580046 363622 580102
rect 363678 580046 381250 580102
rect 381306 580046 381374 580102
rect 381430 580046 381498 580102
rect 381554 580046 381622 580102
rect 381678 580046 399250 580102
rect 399306 580046 399374 580102
rect 399430 580046 399498 580102
rect 399554 580046 399622 580102
rect 399678 580046 417250 580102
rect 417306 580046 417374 580102
rect 417430 580046 417498 580102
rect 417554 580046 417622 580102
rect 417678 580046 435250 580102
rect 435306 580046 435374 580102
rect 435430 580046 435498 580102
rect 435554 580046 435622 580102
rect 435678 580046 453250 580102
rect 453306 580046 453374 580102
rect 453430 580046 453498 580102
rect 453554 580046 453622 580102
rect 453678 580046 471250 580102
rect 471306 580046 471374 580102
rect 471430 580046 471498 580102
rect 471554 580046 471622 580102
rect 471678 580046 489250 580102
rect 489306 580046 489374 580102
rect 489430 580046 489498 580102
rect 489554 580046 489622 580102
rect 489678 580046 507250 580102
rect 507306 580046 507374 580102
rect 507430 580046 507498 580102
rect 507554 580046 507622 580102
rect 507678 580046 525250 580102
rect 525306 580046 525374 580102
rect 525430 580046 525498 580102
rect 525554 580046 525622 580102
rect 525678 580046 543250 580102
rect 543306 580046 543374 580102
rect 543430 580046 543498 580102
rect 543554 580046 543622 580102
rect 543678 580046 561250 580102
rect 561306 580046 561374 580102
rect 561430 580046 561498 580102
rect 561554 580046 561622 580102
rect 561678 580046 579250 580102
rect 579306 580046 579374 580102
rect 579430 580046 579498 580102
rect 579554 580046 579622 580102
rect 579678 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597980 580102
rect -1916 579978 597980 580046
rect -1916 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 3250 579978
rect 3306 579922 3374 579978
rect 3430 579922 3498 579978
rect 3554 579922 3622 579978
rect 3678 579922 21250 579978
rect 21306 579922 21374 579978
rect 21430 579922 21498 579978
rect 21554 579922 21622 579978
rect 21678 579922 39250 579978
rect 39306 579922 39374 579978
rect 39430 579922 39498 579978
rect 39554 579922 39622 579978
rect 39678 579922 57250 579978
rect 57306 579922 57374 579978
rect 57430 579922 57498 579978
rect 57554 579922 57622 579978
rect 57678 579922 75250 579978
rect 75306 579922 75374 579978
rect 75430 579922 75498 579978
rect 75554 579922 75622 579978
rect 75678 579922 93250 579978
rect 93306 579922 93374 579978
rect 93430 579922 93498 579978
rect 93554 579922 93622 579978
rect 93678 579922 111250 579978
rect 111306 579922 111374 579978
rect 111430 579922 111498 579978
rect 111554 579922 111622 579978
rect 111678 579922 129250 579978
rect 129306 579922 129374 579978
rect 129430 579922 129498 579978
rect 129554 579922 129622 579978
rect 129678 579922 147250 579978
rect 147306 579922 147374 579978
rect 147430 579922 147498 579978
rect 147554 579922 147622 579978
rect 147678 579922 165250 579978
rect 165306 579922 165374 579978
rect 165430 579922 165498 579978
rect 165554 579922 165622 579978
rect 165678 579922 183250 579978
rect 183306 579922 183374 579978
rect 183430 579922 183498 579978
rect 183554 579922 183622 579978
rect 183678 579922 201250 579978
rect 201306 579922 201374 579978
rect 201430 579922 201498 579978
rect 201554 579922 201622 579978
rect 201678 579922 219250 579978
rect 219306 579922 219374 579978
rect 219430 579922 219498 579978
rect 219554 579922 219622 579978
rect 219678 579922 237250 579978
rect 237306 579922 237374 579978
rect 237430 579922 237498 579978
rect 237554 579922 237622 579978
rect 237678 579922 255250 579978
rect 255306 579922 255374 579978
rect 255430 579922 255498 579978
rect 255554 579922 255622 579978
rect 255678 579922 273250 579978
rect 273306 579922 273374 579978
rect 273430 579922 273498 579978
rect 273554 579922 273622 579978
rect 273678 579922 291250 579978
rect 291306 579922 291374 579978
rect 291430 579922 291498 579978
rect 291554 579922 291622 579978
rect 291678 579922 309250 579978
rect 309306 579922 309374 579978
rect 309430 579922 309498 579978
rect 309554 579922 309622 579978
rect 309678 579922 327250 579978
rect 327306 579922 327374 579978
rect 327430 579922 327498 579978
rect 327554 579922 327622 579978
rect 327678 579922 345250 579978
rect 345306 579922 345374 579978
rect 345430 579922 345498 579978
rect 345554 579922 345622 579978
rect 345678 579922 363250 579978
rect 363306 579922 363374 579978
rect 363430 579922 363498 579978
rect 363554 579922 363622 579978
rect 363678 579922 381250 579978
rect 381306 579922 381374 579978
rect 381430 579922 381498 579978
rect 381554 579922 381622 579978
rect 381678 579922 399250 579978
rect 399306 579922 399374 579978
rect 399430 579922 399498 579978
rect 399554 579922 399622 579978
rect 399678 579922 417250 579978
rect 417306 579922 417374 579978
rect 417430 579922 417498 579978
rect 417554 579922 417622 579978
rect 417678 579922 435250 579978
rect 435306 579922 435374 579978
rect 435430 579922 435498 579978
rect 435554 579922 435622 579978
rect 435678 579922 453250 579978
rect 453306 579922 453374 579978
rect 453430 579922 453498 579978
rect 453554 579922 453622 579978
rect 453678 579922 471250 579978
rect 471306 579922 471374 579978
rect 471430 579922 471498 579978
rect 471554 579922 471622 579978
rect 471678 579922 489250 579978
rect 489306 579922 489374 579978
rect 489430 579922 489498 579978
rect 489554 579922 489622 579978
rect 489678 579922 507250 579978
rect 507306 579922 507374 579978
rect 507430 579922 507498 579978
rect 507554 579922 507622 579978
rect 507678 579922 525250 579978
rect 525306 579922 525374 579978
rect 525430 579922 525498 579978
rect 525554 579922 525622 579978
rect 525678 579922 543250 579978
rect 543306 579922 543374 579978
rect 543430 579922 543498 579978
rect 543554 579922 543622 579978
rect 543678 579922 561250 579978
rect 561306 579922 561374 579978
rect 561430 579922 561498 579978
rect 561554 579922 561622 579978
rect 561678 579922 579250 579978
rect 579306 579922 579374 579978
rect 579430 579922 579498 579978
rect 579554 579922 579622 579978
rect 579678 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597980 579978
rect -1916 579826 597980 579922
rect -1916 568350 597980 568446
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 6970 568350
rect 7026 568294 7094 568350
rect 7150 568294 7218 568350
rect 7274 568294 7342 568350
rect 7398 568294 24970 568350
rect 25026 568294 25094 568350
rect 25150 568294 25218 568350
rect 25274 568294 25342 568350
rect 25398 568294 42970 568350
rect 43026 568294 43094 568350
rect 43150 568294 43218 568350
rect 43274 568294 43342 568350
rect 43398 568294 60970 568350
rect 61026 568294 61094 568350
rect 61150 568294 61218 568350
rect 61274 568294 61342 568350
rect 61398 568294 78970 568350
rect 79026 568294 79094 568350
rect 79150 568294 79218 568350
rect 79274 568294 79342 568350
rect 79398 568294 96970 568350
rect 97026 568294 97094 568350
rect 97150 568294 97218 568350
rect 97274 568294 97342 568350
rect 97398 568294 114970 568350
rect 115026 568294 115094 568350
rect 115150 568294 115218 568350
rect 115274 568294 115342 568350
rect 115398 568294 132970 568350
rect 133026 568294 133094 568350
rect 133150 568294 133218 568350
rect 133274 568294 133342 568350
rect 133398 568294 150970 568350
rect 151026 568294 151094 568350
rect 151150 568294 151218 568350
rect 151274 568294 151342 568350
rect 151398 568294 168970 568350
rect 169026 568294 169094 568350
rect 169150 568294 169218 568350
rect 169274 568294 169342 568350
rect 169398 568294 186970 568350
rect 187026 568294 187094 568350
rect 187150 568294 187218 568350
rect 187274 568294 187342 568350
rect 187398 568294 204970 568350
rect 205026 568294 205094 568350
rect 205150 568294 205218 568350
rect 205274 568294 205342 568350
rect 205398 568294 222970 568350
rect 223026 568294 223094 568350
rect 223150 568294 223218 568350
rect 223274 568294 223342 568350
rect 223398 568294 240970 568350
rect 241026 568294 241094 568350
rect 241150 568294 241218 568350
rect 241274 568294 241342 568350
rect 241398 568294 258970 568350
rect 259026 568294 259094 568350
rect 259150 568294 259218 568350
rect 259274 568294 259342 568350
rect 259398 568294 276970 568350
rect 277026 568294 277094 568350
rect 277150 568294 277218 568350
rect 277274 568294 277342 568350
rect 277398 568294 294970 568350
rect 295026 568294 295094 568350
rect 295150 568294 295218 568350
rect 295274 568294 295342 568350
rect 295398 568294 312970 568350
rect 313026 568294 313094 568350
rect 313150 568294 313218 568350
rect 313274 568294 313342 568350
rect 313398 568294 330970 568350
rect 331026 568294 331094 568350
rect 331150 568294 331218 568350
rect 331274 568294 331342 568350
rect 331398 568294 348970 568350
rect 349026 568294 349094 568350
rect 349150 568294 349218 568350
rect 349274 568294 349342 568350
rect 349398 568294 366970 568350
rect 367026 568294 367094 568350
rect 367150 568294 367218 568350
rect 367274 568294 367342 568350
rect 367398 568294 384970 568350
rect 385026 568294 385094 568350
rect 385150 568294 385218 568350
rect 385274 568294 385342 568350
rect 385398 568294 402970 568350
rect 403026 568294 403094 568350
rect 403150 568294 403218 568350
rect 403274 568294 403342 568350
rect 403398 568294 420970 568350
rect 421026 568294 421094 568350
rect 421150 568294 421218 568350
rect 421274 568294 421342 568350
rect 421398 568294 438970 568350
rect 439026 568294 439094 568350
rect 439150 568294 439218 568350
rect 439274 568294 439342 568350
rect 439398 568294 456970 568350
rect 457026 568294 457094 568350
rect 457150 568294 457218 568350
rect 457274 568294 457342 568350
rect 457398 568294 474970 568350
rect 475026 568294 475094 568350
rect 475150 568294 475218 568350
rect 475274 568294 475342 568350
rect 475398 568294 492970 568350
rect 493026 568294 493094 568350
rect 493150 568294 493218 568350
rect 493274 568294 493342 568350
rect 493398 568294 510970 568350
rect 511026 568294 511094 568350
rect 511150 568294 511218 568350
rect 511274 568294 511342 568350
rect 511398 568294 528970 568350
rect 529026 568294 529094 568350
rect 529150 568294 529218 568350
rect 529274 568294 529342 568350
rect 529398 568294 546970 568350
rect 547026 568294 547094 568350
rect 547150 568294 547218 568350
rect 547274 568294 547342 568350
rect 547398 568294 564970 568350
rect 565026 568294 565094 568350
rect 565150 568294 565218 568350
rect 565274 568294 565342 568350
rect 565398 568294 582970 568350
rect 583026 568294 583094 568350
rect 583150 568294 583218 568350
rect 583274 568294 583342 568350
rect 583398 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect -1916 568226 597980 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 6970 568226
rect 7026 568170 7094 568226
rect 7150 568170 7218 568226
rect 7274 568170 7342 568226
rect 7398 568170 24970 568226
rect 25026 568170 25094 568226
rect 25150 568170 25218 568226
rect 25274 568170 25342 568226
rect 25398 568170 42970 568226
rect 43026 568170 43094 568226
rect 43150 568170 43218 568226
rect 43274 568170 43342 568226
rect 43398 568170 60970 568226
rect 61026 568170 61094 568226
rect 61150 568170 61218 568226
rect 61274 568170 61342 568226
rect 61398 568170 78970 568226
rect 79026 568170 79094 568226
rect 79150 568170 79218 568226
rect 79274 568170 79342 568226
rect 79398 568170 96970 568226
rect 97026 568170 97094 568226
rect 97150 568170 97218 568226
rect 97274 568170 97342 568226
rect 97398 568170 114970 568226
rect 115026 568170 115094 568226
rect 115150 568170 115218 568226
rect 115274 568170 115342 568226
rect 115398 568170 132970 568226
rect 133026 568170 133094 568226
rect 133150 568170 133218 568226
rect 133274 568170 133342 568226
rect 133398 568170 150970 568226
rect 151026 568170 151094 568226
rect 151150 568170 151218 568226
rect 151274 568170 151342 568226
rect 151398 568170 168970 568226
rect 169026 568170 169094 568226
rect 169150 568170 169218 568226
rect 169274 568170 169342 568226
rect 169398 568170 186970 568226
rect 187026 568170 187094 568226
rect 187150 568170 187218 568226
rect 187274 568170 187342 568226
rect 187398 568170 204970 568226
rect 205026 568170 205094 568226
rect 205150 568170 205218 568226
rect 205274 568170 205342 568226
rect 205398 568170 222970 568226
rect 223026 568170 223094 568226
rect 223150 568170 223218 568226
rect 223274 568170 223342 568226
rect 223398 568170 240970 568226
rect 241026 568170 241094 568226
rect 241150 568170 241218 568226
rect 241274 568170 241342 568226
rect 241398 568170 258970 568226
rect 259026 568170 259094 568226
rect 259150 568170 259218 568226
rect 259274 568170 259342 568226
rect 259398 568170 276970 568226
rect 277026 568170 277094 568226
rect 277150 568170 277218 568226
rect 277274 568170 277342 568226
rect 277398 568170 294970 568226
rect 295026 568170 295094 568226
rect 295150 568170 295218 568226
rect 295274 568170 295342 568226
rect 295398 568170 312970 568226
rect 313026 568170 313094 568226
rect 313150 568170 313218 568226
rect 313274 568170 313342 568226
rect 313398 568170 330970 568226
rect 331026 568170 331094 568226
rect 331150 568170 331218 568226
rect 331274 568170 331342 568226
rect 331398 568170 348970 568226
rect 349026 568170 349094 568226
rect 349150 568170 349218 568226
rect 349274 568170 349342 568226
rect 349398 568170 366970 568226
rect 367026 568170 367094 568226
rect 367150 568170 367218 568226
rect 367274 568170 367342 568226
rect 367398 568170 384970 568226
rect 385026 568170 385094 568226
rect 385150 568170 385218 568226
rect 385274 568170 385342 568226
rect 385398 568170 402970 568226
rect 403026 568170 403094 568226
rect 403150 568170 403218 568226
rect 403274 568170 403342 568226
rect 403398 568170 420970 568226
rect 421026 568170 421094 568226
rect 421150 568170 421218 568226
rect 421274 568170 421342 568226
rect 421398 568170 438970 568226
rect 439026 568170 439094 568226
rect 439150 568170 439218 568226
rect 439274 568170 439342 568226
rect 439398 568170 456970 568226
rect 457026 568170 457094 568226
rect 457150 568170 457218 568226
rect 457274 568170 457342 568226
rect 457398 568170 474970 568226
rect 475026 568170 475094 568226
rect 475150 568170 475218 568226
rect 475274 568170 475342 568226
rect 475398 568170 492970 568226
rect 493026 568170 493094 568226
rect 493150 568170 493218 568226
rect 493274 568170 493342 568226
rect 493398 568170 510970 568226
rect 511026 568170 511094 568226
rect 511150 568170 511218 568226
rect 511274 568170 511342 568226
rect 511398 568170 528970 568226
rect 529026 568170 529094 568226
rect 529150 568170 529218 568226
rect 529274 568170 529342 568226
rect 529398 568170 546970 568226
rect 547026 568170 547094 568226
rect 547150 568170 547218 568226
rect 547274 568170 547342 568226
rect 547398 568170 564970 568226
rect 565026 568170 565094 568226
rect 565150 568170 565218 568226
rect 565274 568170 565342 568226
rect 565398 568170 582970 568226
rect 583026 568170 583094 568226
rect 583150 568170 583218 568226
rect 583274 568170 583342 568226
rect 583398 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect -1916 568102 597980 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 6970 568102
rect 7026 568046 7094 568102
rect 7150 568046 7218 568102
rect 7274 568046 7342 568102
rect 7398 568046 24970 568102
rect 25026 568046 25094 568102
rect 25150 568046 25218 568102
rect 25274 568046 25342 568102
rect 25398 568046 42970 568102
rect 43026 568046 43094 568102
rect 43150 568046 43218 568102
rect 43274 568046 43342 568102
rect 43398 568046 60970 568102
rect 61026 568046 61094 568102
rect 61150 568046 61218 568102
rect 61274 568046 61342 568102
rect 61398 568046 78970 568102
rect 79026 568046 79094 568102
rect 79150 568046 79218 568102
rect 79274 568046 79342 568102
rect 79398 568046 96970 568102
rect 97026 568046 97094 568102
rect 97150 568046 97218 568102
rect 97274 568046 97342 568102
rect 97398 568046 114970 568102
rect 115026 568046 115094 568102
rect 115150 568046 115218 568102
rect 115274 568046 115342 568102
rect 115398 568046 132970 568102
rect 133026 568046 133094 568102
rect 133150 568046 133218 568102
rect 133274 568046 133342 568102
rect 133398 568046 150970 568102
rect 151026 568046 151094 568102
rect 151150 568046 151218 568102
rect 151274 568046 151342 568102
rect 151398 568046 168970 568102
rect 169026 568046 169094 568102
rect 169150 568046 169218 568102
rect 169274 568046 169342 568102
rect 169398 568046 186970 568102
rect 187026 568046 187094 568102
rect 187150 568046 187218 568102
rect 187274 568046 187342 568102
rect 187398 568046 204970 568102
rect 205026 568046 205094 568102
rect 205150 568046 205218 568102
rect 205274 568046 205342 568102
rect 205398 568046 222970 568102
rect 223026 568046 223094 568102
rect 223150 568046 223218 568102
rect 223274 568046 223342 568102
rect 223398 568046 240970 568102
rect 241026 568046 241094 568102
rect 241150 568046 241218 568102
rect 241274 568046 241342 568102
rect 241398 568046 258970 568102
rect 259026 568046 259094 568102
rect 259150 568046 259218 568102
rect 259274 568046 259342 568102
rect 259398 568046 276970 568102
rect 277026 568046 277094 568102
rect 277150 568046 277218 568102
rect 277274 568046 277342 568102
rect 277398 568046 294970 568102
rect 295026 568046 295094 568102
rect 295150 568046 295218 568102
rect 295274 568046 295342 568102
rect 295398 568046 312970 568102
rect 313026 568046 313094 568102
rect 313150 568046 313218 568102
rect 313274 568046 313342 568102
rect 313398 568046 330970 568102
rect 331026 568046 331094 568102
rect 331150 568046 331218 568102
rect 331274 568046 331342 568102
rect 331398 568046 348970 568102
rect 349026 568046 349094 568102
rect 349150 568046 349218 568102
rect 349274 568046 349342 568102
rect 349398 568046 366970 568102
rect 367026 568046 367094 568102
rect 367150 568046 367218 568102
rect 367274 568046 367342 568102
rect 367398 568046 384970 568102
rect 385026 568046 385094 568102
rect 385150 568046 385218 568102
rect 385274 568046 385342 568102
rect 385398 568046 402970 568102
rect 403026 568046 403094 568102
rect 403150 568046 403218 568102
rect 403274 568046 403342 568102
rect 403398 568046 420970 568102
rect 421026 568046 421094 568102
rect 421150 568046 421218 568102
rect 421274 568046 421342 568102
rect 421398 568046 438970 568102
rect 439026 568046 439094 568102
rect 439150 568046 439218 568102
rect 439274 568046 439342 568102
rect 439398 568046 456970 568102
rect 457026 568046 457094 568102
rect 457150 568046 457218 568102
rect 457274 568046 457342 568102
rect 457398 568046 474970 568102
rect 475026 568046 475094 568102
rect 475150 568046 475218 568102
rect 475274 568046 475342 568102
rect 475398 568046 492970 568102
rect 493026 568046 493094 568102
rect 493150 568046 493218 568102
rect 493274 568046 493342 568102
rect 493398 568046 510970 568102
rect 511026 568046 511094 568102
rect 511150 568046 511218 568102
rect 511274 568046 511342 568102
rect 511398 568046 528970 568102
rect 529026 568046 529094 568102
rect 529150 568046 529218 568102
rect 529274 568046 529342 568102
rect 529398 568046 546970 568102
rect 547026 568046 547094 568102
rect 547150 568046 547218 568102
rect 547274 568046 547342 568102
rect 547398 568046 564970 568102
rect 565026 568046 565094 568102
rect 565150 568046 565218 568102
rect 565274 568046 565342 568102
rect 565398 568046 582970 568102
rect 583026 568046 583094 568102
rect 583150 568046 583218 568102
rect 583274 568046 583342 568102
rect 583398 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect -1916 567978 597980 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 6970 567978
rect 7026 567922 7094 567978
rect 7150 567922 7218 567978
rect 7274 567922 7342 567978
rect 7398 567922 24970 567978
rect 25026 567922 25094 567978
rect 25150 567922 25218 567978
rect 25274 567922 25342 567978
rect 25398 567922 42970 567978
rect 43026 567922 43094 567978
rect 43150 567922 43218 567978
rect 43274 567922 43342 567978
rect 43398 567922 60970 567978
rect 61026 567922 61094 567978
rect 61150 567922 61218 567978
rect 61274 567922 61342 567978
rect 61398 567922 78970 567978
rect 79026 567922 79094 567978
rect 79150 567922 79218 567978
rect 79274 567922 79342 567978
rect 79398 567922 96970 567978
rect 97026 567922 97094 567978
rect 97150 567922 97218 567978
rect 97274 567922 97342 567978
rect 97398 567922 114970 567978
rect 115026 567922 115094 567978
rect 115150 567922 115218 567978
rect 115274 567922 115342 567978
rect 115398 567922 132970 567978
rect 133026 567922 133094 567978
rect 133150 567922 133218 567978
rect 133274 567922 133342 567978
rect 133398 567922 150970 567978
rect 151026 567922 151094 567978
rect 151150 567922 151218 567978
rect 151274 567922 151342 567978
rect 151398 567922 168970 567978
rect 169026 567922 169094 567978
rect 169150 567922 169218 567978
rect 169274 567922 169342 567978
rect 169398 567922 186970 567978
rect 187026 567922 187094 567978
rect 187150 567922 187218 567978
rect 187274 567922 187342 567978
rect 187398 567922 204970 567978
rect 205026 567922 205094 567978
rect 205150 567922 205218 567978
rect 205274 567922 205342 567978
rect 205398 567922 222970 567978
rect 223026 567922 223094 567978
rect 223150 567922 223218 567978
rect 223274 567922 223342 567978
rect 223398 567922 240970 567978
rect 241026 567922 241094 567978
rect 241150 567922 241218 567978
rect 241274 567922 241342 567978
rect 241398 567922 258970 567978
rect 259026 567922 259094 567978
rect 259150 567922 259218 567978
rect 259274 567922 259342 567978
rect 259398 567922 276970 567978
rect 277026 567922 277094 567978
rect 277150 567922 277218 567978
rect 277274 567922 277342 567978
rect 277398 567922 294970 567978
rect 295026 567922 295094 567978
rect 295150 567922 295218 567978
rect 295274 567922 295342 567978
rect 295398 567922 312970 567978
rect 313026 567922 313094 567978
rect 313150 567922 313218 567978
rect 313274 567922 313342 567978
rect 313398 567922 330970 567978
rect 331026 567922 331094 567978
rect 331150 567922 331218 567978
rect 331274 567922 331342 567978
rect 331398 567922 348970 567978
rect 349026 567922 349094 567978
rect 349150 567922 349218 567978
rect 349274 567922 349342 567978
rect 349398 567922 366970 567978
rect 367026 567922 367094 567978
rect 367150 567922 367218 567978
rect 367274 567922 367342 567978
rect 367398 567922 384970 567978
rect 385026 567922 385094 567978
rect 385150 567922 385218 567978
rect 385274 567922 385342 567978
rect 385398 567922 402970 567978
rect 403026 567922 403094 567978
rect 403150 567922 403218 567978
rect 403274 567922 403342 567978
rect 403398 567922 420970 567978
rect 421026 567922 421094 567978
rect 421150 567922 421218 567978
rect 421274 567922 421342 567978
rect 421398 567922 438970 567978
rect 439026 567922 439094 567978
rect 439150 567922 439218 567978
rect 439274 567922 439342 567978
rect 439398 567922 456970 567978
rect 457026 567922 457094 567978
rect 457150 567922 457218 567978
rect 457274 567922 457342 567978
rect 457398 567922 474970 567978
rect 475026 567922 475094 567978
rect 475150 567922 475218 567978
rect 475274 567922 475342 567978
rect 475398 567922 492970 567978
rect 493026 567922 493094 567978
rect 493150 567922 493218 567978
rect 493274 567922 493342 567978
rect 493398 567922 510970 567978
rect 511026 567922 511094 567978
rect 511150 567922 511218 567978
rect 511274 567922 511342 567978
rect 511398 567922 528970 567978
rect 529026 567922 529094 567978
rect 529150 567922 529218 567978
rect 529274 567922 529342 567978
rect 529398 567922 546970 567978
rect 547026 567922 547094 567978
rect 547150 567922 547218 567978
rect 547274 567922 547342 567978
rect 547398 567922 564970 567978
rect 565026 567922 565094 567978
rect 565150 567922 565218 567978
rect 565274 567922 565342 567978
rect 565398 567922 582970 567978
rect 583026 567922 583094 567978
rect 583150 567922 583218 567978
rect 583274 567922 583342 567978
rect 583398 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect -1916 567826 597980 567922
rect -1916 562350 597980 562446
rect -1916 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 3250 562350
rect 3306 562294 3374 562350
rect 3430 562294 3498 562350
rect 3554 562294 3622 562350
rect 3678 562294 21250 562350
rect 21306 562294 21374 562350
rect 21430 562294 21498 562350
rect 21554 562294 21622 562350
rect 21678 562294 39250 562350
rect 39306 562294 39374 562350
rect 39430 562294 39498 562350
rect 39554 562294 39622 562350
rect 39678 562294 57250 562350
rect 57306 562294 57374 562350
rect 57430 562294 57498 562350
rect 57554 562294 57622 562350
rect 57678 562294 75250 562350
rect 75306 562294 75374 562350
rect 75430 562294 75498 562350
rect 75554 562294 75622 562350
rect 75678 562294 93250 562350
rect 93306 562294 93374 562350
rect 93430 562294 93498 562350
rect 93554 562294 93622 562350
rect 93678 562294 111250 562350
rect 111306 562294 111374 562350
rect 111430 562294 111498 562350
rect 111554 562294 111622 562350
rect 111678 562294 129250 562350
rect 129306 562294 129374 562350
rect 129430 562294 129498 562350
rect 129554 562294 129622 562350
rect 129678 562294 147250 562350
rect 147306 562294 147374 562350
rect 147430 562294 147498 562350
rect 147554 562294 147622 562350
rect 147678 562294 165250 562350
rect 165306 562294 165374 562350
rect 165430 562294 165498 562350
rect 165554 562294 165622 562350
rect 165678 562294 183250 562350
rect 183306 562294 183374 562350
rect 183430 562294 183498 562350
rect 183554 562294 183622 562350
rect 183678 562294 201250 562350
rect 201306 562294 201374 562350
rect 201430 562294 201498 562350
rect 201554 562294 201622 562350
rect 201678 562294 219250 562350
rect 219306 562294 219374 562350
rect 219430 562294 219498 562350
rect 219554 562294 219622 562350
rect 219678 562294 237250 562350
rect 237306 562294 237374 562350
rect 237430 562294 237498 562350
rect 237554 562294 237622 562350
rect 237678 562294 255250 562350
rect 255306 562294 255374 562350
rect 255430 562294 255498 562350
rect 255554 562294 255622 562350
rect 255678 562294 273250 562350
rect 273306 562294 273374 562350
rect 273430 562294 273498 562350
rect 273554 562294 273622 562350
rect 273678 562294 291250 562350
rect 291306 562294 291374 562350
rect 291430 562294 291498 562350
rect 291554 562294 291622 562350
rect 291678 562294 309250 562350
rect 309306 562294 309374 562350
rect 309430 562294 309498 562350
rect 309554 562294 309622 562350
rect 309678 562294 327250 562350
rect 327306 562294 327374 562350
rect 327430 562294 327498 562350
rect 327554 562294 327622 562350
rect 327678 562294 345250 562350
rect 345306 562294 345374 562350
rect 345430 562294 345498 562350
rect 345554 562294 345622 562350
rect 345678 562294 363250 562350
rect 363306 562294 363374 562350
rect 363430 562294 363498 562350
rect 363554 562294 363622 562350
rect 363678 562294 381250 562350
rect 381306 562294 381374 562350
rect 381430 562294 381498 562350
rect 381554 562294 381622 562350
rect 381678 562294 399250 562350
rect 399306 562294 399374 562350
rect 399430 562294 399498 562350
rect 399554 562294 399622 562350
rect 399678 562294 417250 562350
rect 417306 562294 417374 562350
rect 417430 562294 417498 562350
rect 417554 562294 417622 562350
rect 417678 562294 435250 562350
rect 435306 562294 435374 562350
rect 435430 562294 435498 562350
rect 435554 562294 435622 562350
rect 435678 562294 453250 562350
rect 453306 562294 453374 562350
rect 453430 562294 453498 562350
rect 453554 562294 453622 562350
rect 453678 562294 471250 562350
rect 471306 562294 471374 562350
rect 471430 562294 471498 562350
rect 471554 562294 471622 562350
rect 471678 562294 489250 562350
rect 489306 562294 489374 562350
rect 489430 562294 489498 562350
rect 489554 562294 489622 562350
rect 489678 562294 507250 562350
rect 507306 562294 507374 562350
rect 507430 562294 507498 562350
rect 507554 562294 507622 562350
rect 507678 562294 525250 562350
rect 525306 562294 525374 562350
rect 525430 562294 525498 562350
rect 525554 562294 525622 562350
rect 525678 562294 543250 562350
rect 543306 562294 543374 562350
rect 543430 562294 543498 562350
rect 543554 562294 543622 562350
rect 543678 562294 561250 562350
rect 561306 562294 561374 562350
rect 561430 562294 561498 562350
rect 561554 562294 561622 562350
rect 561678 562294 579250 562350
rect 579306 562294 579374 562350
rect 579430 562294 579498 562350
rect 579554 562294 579622 562350
rect 579678 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597980 562350
rect -1916 562226 597980 562294
rect -1916 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 3250 562226
rect 3306 562170 3374 562226
rect 3430 562170 3498 562226
rect 3554 562170 3622 562226
rect 3678 562170 21250 562226
rect 21306 562170 21374 562226
rect 21430 562170 21498 562226
rect 21554 562170 21622 562226
rect 21678 562170 39250 562226
rect 39306 562170 39374 562226
rect 39430 562170 39498 562226
rect 39554 562170 39622 562226
rect 39678 562170 57250 562226
rect 57306 562170 57374 562226
rect 57430 562170 57498 562226
rect 57554 562170 57622 562226
rect 57678 562170 75250 562226
rect 75306 562170 75374 562226
rect 75430 562170 75498 562226
rect 75554 562170 75622 562226
rect 75678 562170 93250 562226
rect 93306 562170 93374 562226
rect 93430 562170 93498 562226
rect 93554 562170 93622 562226
rect 93678 562170 111250 562226
rect 111306 562170 111374 562226
rect 111430 562170 111498 562226
rect 111554 562170 111622 562226
rect 111678 562170 129250 562226
rect 129306 562170 129374 562226
rect 129430 562170 129498 562226
rect 129554 562170 129622 562226
rect 129678 562170 147250 562226
rect 147306 562170 147374 562226
rect 147430 562170 147498 562226
rect 147554 562170 147622 562226
rect 147678 562170 165250 562226
rect 165306 562170 165374 562226
rect 165430 562170 165498 562226
rect 165554 562170 165622 562226
rect 165678 562170 183250 562226
rect 183306 562170 183374 562226
rect 183430 562170 183498 562226
rect 183554 562170 183622 562226
rect 183678 562170 201250 562226
rect 201306 562170 201374 562226
rect 201430 562170 201498 562226
rect 201554 562170 201622 562226
rect 201678 562170 219250 562226
rect 219306 562170 219374 562226
rect 219430 562170 219498 562226
rect 219554 562170 219622 562226
rect 219678 562170 237250 562226
rect 237306 562170 237374 562226
rect 237430 562170 237498 562226
rect 237554 562170 237622 562226
rect 237678 562170 255250 562226
rect 255306 562170 255374 562226
rect 255430 562170 255498 562226
rect 255554 562170 255622 562226
rect 255678 562170 273250 562226
rect 273306 562170 273374 562226
rect 273430 562170 273498 562226
rect 273554 562170 273622 562226
rect 273678 562170 291250 562226
rect 291306 562170 291374 562226
rect 291430 562170 291498 562226
rect 291554 562170 291622 562226
rect 291678 562170 309250 562226
rect 309306 562170 309374 562226
rect 309430 562170 309498 562226
rect 309554 562170 309622 562226
rect 309678 562170 327250 562226
rect 327306 562170 327374 562226
rect 327430 562170 327498 562226
rect 327554 562170 327622 562226
rect 327678 562170 345250 562226
rect 345306 562170 345374 562226
rect 345430 562170 345498 562226
rect 345554 562170 345622 562226
rect 345678 562170 363250 562226
rect 363306 562170 363374 562226
rect 363430 562170 363498 562226
rect 363554 562170 363622 562226
rect 363678 562170 381250 562226
rect 381306 562170 381374 562226
rect 381430 562170 381498 562226
rect 381554 562170 381622 562226
rect 381678 562170 399250 562226
rect 399306 562170 399374 562226
rect 399430 562170 399498 562226
rect 399554 562170 399622 562226
rect 399678 562170 417250 562226
rect 417306 562170 417374 562226
rect 417430 562170 417498 562226
rect 417554 562170 417622 562226
rect 417678 562170 435250 562226
rect 435306 562170 435374 562226
rect 435430 562170 435498 562226
rect 435554 562170 435622 562226
rect 435678 562170 453250 562226
rect 453306 562170 453374 562226
rect 453430 562170 453498 562226
rect 453554 562170 453622 562226
rect 453678 562170 471250 562226
rect 471306 562170 471374 562226
rect 471430 562170 471498 562226
rect 471554 562170 471622 562226
rect 471678 562170 489250 562226
rect 489306 562170 489374 562226
rect 489430 562170 489498 562226
rect 489554 562170 489622 562226
rect 489678 562170 507250 562226
rect 507306 562170 507374 562226
rect 507430 562170 507498 562226
rect 507554 562170 507622 562226
rect 507678 562170 525250 562226
rect 525306 562170 525374 562226
rect 525430 562170 525498 562226
rect 525554 562170 525622 562226
rect 525678 562170 543250 562226
rect 543306 562170 543374 562226
rect 543430 562170 543498 562226
rect 543554 562170 543622 562226
rect 543678 562170 561250 562226
rect 561306 562170 561374 562226
rect 561430 562170 561498 562226
rect 561554 562170 561622 562226
rect 561678 562170 579250 562226
rect 579306 562170 579374 562226
rect 579430 562170 579498 562226
rect 579554 562170 579622 562226
rect 579678 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597980 562226
rect -1916 562102 597980 562170
rect -1916 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 3250 562102
rect 3306 562046 3374 562102
rect 3430 562046 3498 562102
rect 3554 562046 3622 562102
rect 3678 562046 21250 562102
rect 21306 562046 21374 562102
rect 21430 562046 21498 562102
rect 21554 562046 21622 562102
rect 21678 562046 39250 562102
rect 39306 562046 39374 562102
rect 39430 562046 39498 562102
rect 39554 562046 39622 562102
rect 39678 562046 57250 562102
rect 57306 562046 57374 562102
rect 57430 562046 57498 562102
rect 57554 562046 57622 562102
rect 57678 562046 75250 562102
rect 75306 562046 75374 562102
rect 75430 562046 75498 562102
rect 75554 562046 75622 562102
rect 75678 562046 93250 562102
rect 93306 562046 93374 562102
rect 93430 562046 93498 562102
rect 93554 562046 93622 562102
rect 93678 562046 111250 562102
rect 111306 562046 111374 562102
rect 111430 562046 111498 562102
rect 111554 562046 111622 562102
rect 111678 562046 129250 562102
rect 129306 562046 129374 562102
rect 129430 562046 129498 562102
rect 129554 562046 129622 562102
rect 129678 562046 147250 562102
rect 147306 562046 147374 562102
rect 147430 562046 147498 562102
rect 147554 562046 147622 562102
rect 147678 562046 165250 562102
rect 165306 562046 165374 562102
rect 165430 562046 165498 562102
rect 165554 562046 165622 562102
rect 165678 562046 183250 562102
rect 183306 562046 183374 562102
rect 183430 562046 183498 562102
rect 183554 562046 183622 562102
rect 183678 562046 201250 562102
rect 201306 562046 201374 562102
rect 201430 562046 201498 562102
rect 201554 562046 201622 562102
rect 201678 562046 219250 562102
rect 219306 562046 219374 562102
rect 219430 562046 219498 562102
rect 219554 562046 219622 562102
rect 219678 562046 237250 562102
rect 237306 562046 237374 562102
rect 237430 562046 237498 562102
rect 237554 562046 237622 562102
rect 237678 562046 255250 562102
rect 255306 562046 255374 562102
rect 255430 562046 255498 562102
rect 255554 562046 255622 562102
rect 255678 562046 273250 562102
rect 273306 562046 273374 562102
rect 273430 562046 273498 562102
rect 273554 562046 273622 562102
rect 273678 562046 291250 562102
rect 291306 562046 291374 562102
rect 291430 562046 291498 562102
rect 291554 562046 291622 562102
rect 291678 562046 309250 562102
rect 309306 562046 309374 562102
rect 309430 562046 309498 562102
rect 309554 562046 309622 562102
rect 309678 562046 327250 562102
rect 327306 562046 327374 562102
rect 327430 562046 327498 562102
rect 327554 562046 327622 562102
rect 327678 562046 345250 562102
rect 345306 562046 345374 562102
rect 345430 562046 345498 562102
rect 345554 562046 345622 562102
rect 345678 562046 363250 562102
rect 363306 562046 363374 562102
rect 363430 562046 363498 562102
rect 363554 562046 363622 562102
rect 363678 562046 381250 562102
rect 381306 562046 381374 562102
rect 381430 562046 381498 562102
rect 381554 562046 381622 562102
rect 381678 562046 399250 562102
rect 399306 562046 399374 562102
rect 399430 562046 399498 562102
rect 399554 562046 399622 562102
rect 399678 562046 417250 562102
rect 417306 562046 417374 562102
rect 417430 562046 417498 562102
rect 417554 562046 417622 562102
rect 417678 562046 435250 562102
rect 435306 562046 435374 562102
rect 435430 562046 435498 562102
rect 435554 562046 435622 562102
rect 435678 562046 453250 562102
rect 453306 562046 453374 562102
rect 453430 562046 453498 562102
rect 453554 562046 453622 562102
rect 453678 562046 471250 562102
rect 471306 562046 471374 562102
rect 471430 562046 471498 562102
rect 471554 562046 471622 562102
rect 471678 562046 489250 562102
rect 489306 562046 489374 562102
rect 489430 562046 489498 562102
rect 489554 562046 489622 562102
rect 489678 562046 507250 562102
rect 507306 562046 507374 562102
rect 507430 562046 507498 562102
rect 507554 562046 507622 562102
rect 507678 562046 525250 562102
rect 525306 562046 525374 562102
rect 525430 562046 525498 562102
rect 525554 562046 525622 562102
rect 525678 562046 543250 562102
rect 543306 562046 543374 562102
rect 543430 562046 543498 562102
rect 543554 562046 543622 562102
rect 543678 562046 561250 562102
rect 561306 562046 561374 562102
rect 561430 562046 561498 562102
rect 561554 562046 561622 562102
rect 561678 562046 579250 562102
rect 579306 562046 579374 562102
rect 579430 562046 579498 562102
rect 579554 562046 579622 562102
rect 579678 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597980 562102
rect -1916 561978 597980 562046
rect -1916 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 3250 561978
rect 3306 561922 3374 561978
rect 3430 561922 3498 561978
rect 3554 561922 3622 561978
rect 3678 561922 21250 561978
rect 21306 561922 21374 561978
rect 21430 561922 21498 561978
rect 21554 561922 21622 561978
rect 21678 561922 39250 561978
rect 39306 561922 39374 561978
rect 39430 561922 39498 561978
rect 39554 561922 39622 561978
rect 39678 561922 57250 561978
rect 57306 561922 57374 561978
rect 57430 561922 57498 561978
rect 57554 561922 57622 561978
rect 57678 561922 75250 561978
rect 75306 561922 75374 561978
rect 75430 561922 75498 561978
rect 75554 561922 75622 561978
rect 75678 561922 93250 561978
rect 93306 561922 93374 561978
rect 93430 561922 93498 561978
rect 93554 561922 93622 561978
rect 93678 561922 111250 561978
rect 111306 561922 111374 561978
rect 111430 561922 111498 561978
rect 111554 561922 111622 561978
rect 111678 561922 129250 561978
rect 129306 561922 129374 561978
rect 129430 561922 129498 561978
rect 129554 561922 129622 561978
rect 129678 561922 147250 561978
rect 147306 561922 147374 561978
rect 147430 561922 147498 561978
rect 147554 561922 147622 561978
rect 147678 561922 165250 561978
rect 165306 561922 165374 561978
rect 165430 561922 165498 561978
rect 165554 561922 165622 561978
rect 165678 561922 183250 561978
rect 183306 561922 183374 561978
rect 183430 561922 183498 561978
rect 183554 561922 183622 561978
rect 183678 561922 201250 561978
rect 201306 561922 201374 561978
rect 201430 561922 201498 561978
rect 201554 561922 201622 561978
rect 201678 561922 219250 561978
rect 219306 561922 219374 561978
rect 219430 561922 219498 561978
rect 219554 561922 219622 561978
rect 219678 561922 237250 561978
rect 237306 561922 237374 561978
rect 237430 561922 237498 561978
rect 237554 561922 237622 561978
rect 237678 561922 255250 561978
rect 255306 561922 255374 561978
rect 255430 561922 255498 561978
rect 255554 561922 255622 561978
rect 255678 561922 273250 561978
rect 273306 561922 273374 561978
rect 273430 561922 273498 561978
rect 273554 561922 273622 561978
rect 273678 561922 291250 561978
rect 291306 561922 291374 561978
rect 291430 561922 291498 561978
rect 291554 561922 291622 561978
rect 291678 561922 309250 561978
rect 309306 561922 309374 561978
rect 309430 561922 309498 561978
rect 309554 561922 309622 561978
rect 309678 561922 327250 561978
rect 327306 561922 327374 561978
rect 327430 561922 327498 561978
rect 327554 561922 327622 561978
rect 327678 561922 345250 561978
rect 345306 561922 345374 561978
rect 345430 561922 345498 561978
rect 345554 561922 345622 561978
rect 345678 561922 363250 561978
rect 363306 561922 363374 561978
rect 363430 561922 363498 561978
rect 363554 561922 363622 561978
rect 363678 561922 381250 561978
rect 381306 561922 381374 561978
rect 381430 561922 381498 561978
rect 381554 561922 381622 561978
rect 381678 561922 399250 561978
rect 399306 561922 399374 561978
rect 399430 561922 399498 561978
rect 399554 561922 399622 561978
rect 399678 561922 417250 561978
rect 417306 561922 417374 561978
rect 417430 561922 417498 561978
rect 417554 561922 417622 561978
rect 417678 561922 435250 561978
rect 435306 561922 435374 561978
rect 435430 561922 435498 561978
rect 435554 561922 435622 561978
rect 435678 561922 453250 561978
rect 453306 561922 453374 561978
rect 453430 561922 453498 561978
rect 453554 561922 453622 561978
rect 453678 561922 471250 561978
rect 471306 561922 471374 561978
rect 471430 561922 471498 561978
rect 471554 561922 471622 561978
rect 471678 561922 489250 561978
rect 489306 561922 489374 561978
rect 489430 561922 489498 561978
rect 489554 561922 489622 561978
rect 489678 561922 507250 561978
rect 507306 561922 507374 561978
rect 507430 561922 507498 561978
rect 507554 561922 507622 561978
rect 507678 561922 525250 561978
rect 525306 561922 525374 561978
rect 525430 561922 525498 561978
rect 525554 561922 525622 561978
rect 525678 561922 543250 561978
rect 543306 561922 543374 561978
rect 543430 561922 543498 561978
rect 543554 561922 543622 561978
rect 543678 561922 561250 561978
rect 561306 561922 561374 561978
rect 561430 561922 561498 561978
rect 561554 561922 561622 561978
rect 561678 561922 579250 561978
rect 579306 561922 579374 561978
rect 579430 561922 579498 561978
rect 579554 561922 579622 561978
rect 579678 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597980 561978
rect -1916 561826 597980 561922
rect -1916 550350 597980 550446
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 6970 550350
rect 7026 550294 7094 550350
rect 7150 550294 7218 550350
rect 7274 550294 7342 550350
rect 7398 550294 24970 550350
rect 25026 550294 25094 550350
rect 25150 550294 25218 550350
rect 25274 550294 25342 550350
rect 25398 550294 42970 550350
rect 43026 550294 43094 550350
rect 43150 550294 43218 550350
rect 43274 550294 43342 550350
rect 43398 550294 60970 550350
rect 61026 550294 61094 550350
rect 61150 550294 61218 550350
rect 61274 550294 61342 550350
rect 61398 550294 78970 550350
rect 79026 550294 79094 550350
rect 79150 550294 79218 550350
rect 79274 550294 79342 550350
rect 79398 550294 96970 550350
rect 97026 550294 97094 550350
rect 97150 550294 97218 550350
rect 97274 550294 97342 550350
rect 97398 550294 114970 550350
rect 115026 550294 115094 550350
rect 115150 550294 115218 550350
rect 115274 550294 115342 550350
rect 115398 550294 132970 550350
rect 133026 550294 133094 550350
rect 133150 550294 133218 550350
rect 133274 550294 133342 550350
rect 133398 550294 150970 550350
rect 151026 550294 151094 550350
rect 151150 550294 151218 550350
rect 151274 550294 151342 550350
rect 151398 550294 168970 550350
rect 169026 550294 169094 550350
rect 169150 550294 169218 550350
rect 169274 550294 169342 550350
rect 169398 550294 186970 550350
rect 187026 550294 187094 550350
rect 187150 550294 187218 550350
rect 187274 550294 187342 550350
rect 187398 550294 204970 550350
rect 205026 550294 205094 550350
rect 205150 550294 205218 550350
rect 205274 550294 205342 550350
rect 205398 550294 222970 550350
rect 223026 550294 223094 550350
rect 223150 550294 223218 550350
rect 223274 550294 223342 550350
rect 223398 550294 240970 550350
rect 241026 550294 241094 550350
rect 241150 550294 241218 550350
rect 241274 550294 241342 550350
rect 241398 550294 258970 550350
rect 259026 550294 259094 550350
rect 259150 550294 259218 550350
rect 259274 550294 259342 550350
rect 259398 550294 276970 550350
rect 277026 550294 277094 550350
rect 277150 550294 277218 550350
rect 277274 550294 277342 550350
rect 277398 550294 294970 550350
rect 295026 550294 295094 550350
rect 295150 550294 295218 550350
rect 295274 550294 295342 550350
rect 295398 550294 312970 550350
rect 313026 550294 313094 550350
rect 313150 550294 313218 550350
rect 313274 550294 313342 550350
rect 313398 550294 330970 550350
rect 331026 550294 331094 550350
rect 331150 550294 331218 550350
rect 331274 550294 331342 550350
rect 331398 550294 348970 550350
rect 349026 550294 349094 550350
rect 349150 550294 349218 550350
rect 349274 550294 349342 550350
rect 349398 550294 366970 550350
rect 367026 550294 367094 550350
rect 367150 550294 367218 550350
rect 367274 550294 367342 550350
rect 367398 550294 384970 550350
rect 385026 550294 385094 550350
rect 385150 550294 385218 550350
rect 385274 550294 385342 550350
rect 385398 550294 402970 550350
rect 403026 550294 403094 550350
rect 403150 550294 403218 550350
rect 403274 550294 403342 550350
rect 403398 550294 420970 550350
rect 421026 550294 421094 550350
rect 421150 550294 421218 550350
rect 421274 550294 421342 550350
rect 421398 550294 438970 550350
rect 439026 550294 439094 550350
rect 439150 550294 439218 550350
rect 439274 550294 439342 550350
rect 439398 550294 456970 550350
rect 457026 550294 457094 550350
rect 457150 550294 457218 550350
rect 457274 550294 457342 550350
rect 457398 550294 474970 550350
rect 475026 550294 475094 550350
rect 475150 550294 475218 550350
rect 475274 550294 475342 550350
rect 475398 550294 492970 550350
rect 493026 550294 493094 550350
rect 493150 550294 493218 550350
rect 493274 550294 493342 550350
rect 493398 550294 510970 550350
rect 511026 550294 511094 550350
rect 511150 550294 511218 550350
rect 511274 550294 511342 550350
rect 511398 550294 528970 550350
rect 529026 550294 529094 550350
rect 529150 550294 529218 550350
rect 529274 550294 529342 550350
rect 529398 550294 546970 550350
rect 547026 550294 547094 550350
rect 547150 550294 547218 550350
rect 547274 550294 547342 550350
rect 547398 550294 564970 550350
rect 565026 550294 565094 550350
rect 565150 550294 565218 550350
rect 565274 550294 565342 550350
rect 565398 550294 582970 550350
rect 583026 550294 583094 550350
rect 583150 550294 583218 550350
rect 583274 550294 583342 550350
rect 583398 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect -1916 550226 597980 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 6970 550226
rect 7026 550170 7094 550226
rect 7150 550170 7218 550226
rect 7274 550170 7342 550226
rect 7398 550170 24970 550226
rect 25026 550170 25094 550226
rect 25150 550170 25218 550226
rect 25274 550170 25342 550226
rect 25398 550170 42970 550226
rect 43026 550170 43094 550226
rect 43150 550170 43218 550226
rect 43274 550170 43342 550226
rect 43398 550170 60970 550226
rect 61026 550170 61094 550226
rect 61150 550170 61218 550226
rect 61274 550170 61342 550226
rect 61398 550170 78970 550226
rect 79026 550170 79094 550226
rect 79150 550170 79218 550226
rect 79274 550170 79342 550226
rect 79398 550170 96970 550226
rect 97026 550170 97094 550226
rect 97150 550170 97218 550226
rect 97274 550170 97342 550226
rect 97398 550170 114970 550226
rect 115026 550170 115094 550226
rect 115150 550170 115218 550226
rect 115274 550170 115342 550226
rect 115398 550170 132970 550226
rect 133026 550170 133094 550226
rect 133150 550170 133218 550226
rect 133274 550170 133342 550226
rect 133398 550170 150970 550226
rect 151026 550170 151094 550226
rect 151150 550170 151218 550226
rect 151274 550170 151342 550226
rect 151398 550170 168970 550226
rect 169026 550170 169094 550226
rect 169150 550170 169218 550226
rect 169274 550170 169342 550226
rect 169398 550170 186970 550226
rect 187026 550170 187094 550226
rect 187150 550170 187218 550226
rect 187274 550170 187342 550226
rect 187398 550170 204970 550226
rect 205026 550170 205094 550226
rect 205150 550170 205218 550226
rect 205274 550170 205342 550226
rect 205398 550170 222970 550226
rect 223026 550170 223094 550226
rect 223150 550170 223218 550226
rect 223274 550170 223342 550226
rect 223398 550170 240970 550226
rect 241026 550170 241094 550226
rect 241150 550170 241218 550226
rect 241274 550170 241342 550226
rect 241398 550170 258970 550226
rect 259026 550170 259094 550226
rect 259150 550170 259218 550226
rect 259274 550170 259342 550226
rect 259398 550170 276970 550226
rect 277026 550170 277094 550226
rect 277150 550170 277218 550226
rect 277274 550170 277342 550226
rect 277398 550170 294970 550226
rect 295026 550170 295094 550226
rect 295150 550170 295218 550226
rect 295274 550170 295342 550226
rect 295398 550170 312970 550226
rect 313026 550170 313094 550226
rect 313150 550170 313218 550226
rect 313274 550170 313342 550226
rect 313398 550170 330970 550226
rect 331026 550170 331094 550226
rect 331150 550170 331218 550226
rect 331274 550170 331342 550226
rect 331398 550170 348970 550226
rect 349026 550170 349094 550226
rect 349150 550170 349218 550226
rect 349274 550170 349342 550226
rect 349398 550170 366970 550226
rect 367026 550170 367094 550226
rect 367150 550170 367218 550226
rect 367274 550170 367342 550226
rect 367398 550170 384970 550226
rect 385026 550170 385094 550226
rect 385150 550170 385218 550226
rect 385274 550170 385342 550226
rect 385398 550170 402970 550226
rect 403026 550170 403094 550226
rect 403150 550170 403218 550226
rect 403274 550170 403342 550226
rect 403398 550170 420970 550226
rect 421026 550170 421094 550226
rect 421150 550170 421218 550226
rect 421274 550170 421342 550226
rect 421398 550170 438970 550226
rect 439026 550170 439094 550226
rect 439150 550170 439218 550226
rect 439274 550170 439342 550226
rect 439398 550170 456970 550226
rect 457026 550170 457094 550226
rect 457150 550170 457218 550226
rect 457274 550170 457342 550226
rect 457398 550170 474970 550226
rect 475026 550170 475094 550226
rect 475150 550170 475218 550226
rect 475274 550170 475342 550226
rect 475398 550170 492970 550226
rect 493026 550170 493094 550226
rect 493150 550170 493218 550226
rect 493274 550170 493342 550226
rect 493398 550170 510970 550226
rect 511026 550170 511094 550226
rect 511150 550170 511218 550226
rect 511274 550170 511342 550226
rect 511398 550170 528970 550226
rect 529026 550170 529094 550226
rect 529150 550170 529218 550226
rect 529274 550170 529342 550226
rect 529398 550170 546970 550226
rect 547026 550170 547094 550226
rect 547150 550170 547218 550226
rect 547274 550170 547342 550226
rect 547398 550170 564970 550226
rect 565026 550170 565094 550226
rect 565150 550170 565218 550226
rect 565274 550170 565342 550226
rect 565398 550170 582970 550226
rect 583026 550170 583094 550226
rect 583150 550170 583218 550226
rect 583274 550170 583342 550226
rect 583398 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect -1916 550102 597980 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 6970 550102
rect 7026 550046 7094 550102
rect 7150 550046 7218 550102
rect 7274 550046 7342 550102
rect 7398 550046 24970 550102
rect 25026 550046 25094 550102
rect 25150 550046 25218 550102
rect 25274 550046 25342 550102
rect 25398 550046 42970 550102
rect 43026 550046 43094 550102
rect 43150 550046 43218 550102
rect 43274 550046 43342 550102
rect 43398 550046 60970 550102
rect 61026 550046 61094 550102
rect 61150 550046 61218 550102
rect 61274 550046 61342 550102
rect 61398 550046 78970 550102
rect 79026 550046 79094 550102
rect 79150 550046 79218 550102
rect 79274 550046 79342 550102
rect 79398 550046 96970 550102
rect 97026 550046 97094 550102
rect 97150 550046 97218 550102
rect 97274 550046 97342 550102
rect 97398 550046 114970 550102
rect 115026 550046 115094 550102
rect 115150 550046 115218 550102
rect 115274 550046 115342 550102
rect 115398 550046 132970 550102
rect 133026 550046 133094 550102
rect 133150 550046 133218 550102
rect 133274 550046 133342 550102
rect 133398 550046 150970 550102
rect 151026 550046 151094 550102
rect 151150 550046 151218 550102
rect 151274 550046 151342 550102
rect 151398 550046 168970 550102
rect 169026 550046 169094 550102
rect 169150 550046 169218 550102
rect 169274 550046 169342 550102
rect 169398 550046 186970 550102
rect 187026 550046 187094 550102
rect 187150 550046 187218 550102
rect 187274 550046 187342 550102
rect 187398 550046 204970 550102
rect 205026 550046 205094 550102
rect 205150 550046 205218 550102
rect 205274 550046 205342 550102
rect 205398 550046 222970 550102
rect 223026 550046 223094 550102
rect 223150 550046 223218 550102
rect 223274 550046 223342 550102
rect 223398 550046 240970 550102
rect 241026 550046 241094 550102
rect 241150 550046 241218 550102
rect 241274 550046 241342 550102
rect 241398 550046 258970 550102
rect 259026 550046 259094 550102
rect 259150 550046 259218 550102
rect 259274 550046 259342 550102
rect 259398 550046 276970 550102
rect 277026 550046 277094 550102
rect 277150 550046 277218 550102
rect 277274 550046 277342 550102
rect 277398 550046 294970 550102
rect 295026 550046 295094 550102
rect 295150 550046 295218 550102
rect 295274 550046 295342 550102
rect 295398 550046 312970 550102
rect 313026 550046 313094 550102
rect 313150 550046 313218 550102
rect 313274 550046 313342 550102
rect 313398 550046 330970 550102
rect 331026 550046 331094 550102
rect 331150 550046 331218 550102
rect 331274 550046 331342 550102
rect 331398 550046 348970 550102
rect 349026 550046 349094 550102
rect 349150 550046 349218 550102
rect 349274 550046 349342 550102
rect 349398 550046 366970 550102
rect 367026 550046 367094 550102
rect 367150 550046 367218 550102
rect 367274 550046 367342 550102
rect 367398 550046 384970 550102
rect 385026 550046 385094 550102
rect 385150 550046 385218 550102
rect 385274 550046 385342 550102
rect 385398 550046 402970 550102
rect 403026 550046 403094 550102
rect 403150 550046 403218 550102
rect 403274 550046 403342 550102
rect 403398 550046 420970 550102
rect 421026 550046 421094 550102
rect 421150 550046 421218 550102
rect 421274 550046 421342 550102
rect 421398 550046 438970 550102
rect 439026 550046 439094 550102
rect 439150 550046 439218 550102
rect 439274 550046 439342 550102
rect 439398 550046 456970 550102
rect 457026 550046 457094 550102
rect 457150 550046 457218 550102
rect 457274 550046 457342 550102
rect 457398 550046 474970 550102
rect 475026 550046 475094 550102
rect 475150 550046 475218 550102
rect 475274 550046 475342 550102
rect 475398 550046 492970 550102
rect 493026 550046 493094 550102
rect 493150 550046 493218 550102
rect 493274 550046 493342 550102
rect 493398 550046 510970 550102
rect 511026 550046 511094 550102
rect 511150 550046 511218 550102
rect 511274 550046 511342 550102
rect 511398 550046 528970 550102
rect 529026 550046 529094 550102
rect 529150 550046 529218 550102
rect 529274 550046 529342 550102
rect 529398 550046 546970 550102
rect 547026 550046 547094 550102
rect 547150 550046 547218 550102
rect 547274 550046 547342 550102
rect 547398 550046 564970 550102
rect 565026 550046 565094 550102
rect 565150 550046 565218 550102
rect 565274 550046 565342 550102
rect 565398 550046 582970 550102
rect 583026 550046 583094 550102
rect 583150 550046 583218 550102
rect 583274 550046 583342 550102
rect 583398 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect -1916 549978 597980 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 6970 549978
rect 7026 549922 7094 549978
rect 7150 549922 7218 549978
rect 7274 549922 7342 549978
rect 7398 549922 24970 549978
rect 25026 549922 25094 549978
rect 25150 549922 25218 549978
rect 25274 549922 25342 549978
rect 25398 549922 42970 549978
rect 43026 549922 43094 549978
rect 43150 549922 43218 549978
rect 43274 549922 43342 549978
rect 43398 549922 60970 549978
rect 61026 549922 61094 549978
rect 61150 549922 61218 549978
rect 61274 549922 61342 549978
rect 61398 549922 78970 549978
rect 79026 549922 79094 549978
rect 79150 549922 79218 549978
rect 79274 549922 79342 549978
rect 79398 549922 96970 549978
rect 97026 549922 97094 549978
rect 97150 549922 97218 549978
rect 97274 549922 97342 549978
rect 97398 549922 114970 549978
rect 115026 549922 115094 549978
rect 115150 549922 115218 549978
rect 115274 549922 115342 549978
rect 115398 549922 132970 549978
rect 133026 549922 133094 549978
rect 133150 549922 133218 549978
rect 133274 549922 133342 549978
rect 133398 549922 150970 549978
rect 151026 549922 151094 549978
rect 151150 549922 151218 549978
rect 151274 549922 151342 549978
rect 151398 549922 168970 549978
rect 169026 549922 169094 549978
rect 169150 549922 169218 549978
rect 169274 549922 169342 549978
rect 169398 549922 186970 549978
rect 187026 549922 187094 549978
rect 187150 549922 187218 549978
rect 187274 549922 187342 549978
rect 187398 549922 204970 549978
rect 205026 549922 205094 549978
rect 205150 549922 205218 549978
rect 205274 549922 205342 549978
rect 205398 549922 222970 549978
rect 223026 549922 223094 549978
rect 223150 549922 223218 549978
rect 223274 549922 223342 549978
rect 223398 549922 240970 549978
rect 241026 549922 241094 549978
rect 241150 549922 241218 549978
rect 241274 549922 241342 549978
rect 241398 549922 258970 549978
rect 259026 549922 259094 549978
rect 259150 549922 259218 549978
rect 259274 549922 259342 549978
rect 259398 549922 276970 549978
rect 277026 549922 277094 549978
rect 277150 549922 277218 549978
rect 277274 549922 277342 549978
rect 277398 549922 294970 549978
rect 295026 549922 295094 549978
rect 295150 549922 295218 549978
rect 295274 549922 295342 549978
rect 295398 549922 312970 549978
rect 313026 549922 313094 549978
rect 313150 549922 313218 549978
rect 313274 549922 313342 549978
rect 313398 549922 330970 549978
rect 331026 549922 331094 549978
rect 331150 549922 331218 549978
rect 331274 549922 331342 549978
rect 331398 549922 348970 549978
rect 349026 549922 349094 549978
rect 349150 549922 349218 549978
rect 349274 549922 349342 549978
rect 349398 549922 366970 549978
rect 367026 549922 367094 549978
rect 367150 549922 367218 549978
rect 367274 549922 367342 549978
rect 367398 549922 384970 549978
rect 385026 549922 385094 549978
rect 385150 549922 385218 549978
rect 385274 549922 385342 549978
rect 385398 549922 402970 549978
rect 403026 549922 403094 549978
rect 403150 549922 403218 549978
rect 403274 549922 403342 549978
rect 403398 549922 420970 549978
rect 421026 549922 421094 549978
rect 421150 549922 421218 549978
rect 421274 549922 421342 549978
rect 421398 549922 438970 549978
rect 439026 549922 439094 549978
rect 439150 549922 439218 549978
rect 439274 549922 439342 549978
rect 439398 549922 456970 549978
rect 457026 549922 457094 549978
rect 457150 549922 457218 549978
rect 457274 549922 457342 549978
rect 457398 549922 474970 549978
rect 475026 549922 475094 549978
rect 475150 549922 475218 549978
rect 475274 549922 475342 549978
rect 475398 549922 492970 549978
rect 493026 549922 493094 549978
rect 493150 549922 493218 549978
rect 493274 549922 493342 549978
rect 493398 549922 510970 549978
rect 511026 549922 511094 549978
rect 511150 549922 511218 549978
rect 511274 549922 511342 549978
rect 511398 549922 528970 549978
rect 529026 549922 529094 549978
rect 529150 549922 529218 549978
rect 529274 549922 529342 549978
rect 529398 549922 546970 549978
rect 547026 549922 547094 549978
rect 547150 549922 547218 549978
rect 547274 549922 547342 549978
rect 547398 549922 564970 549978
rect 565026 549922 565094 549978
rect 565150 549922 565218 549978
rect 565274 549922 565342 549978
rect 565398 549922 582970 549978
rect 583026 549922 583094 549978
rect 583150 549922 583218 549978
rect 583274 549922 583342 549978
rect 583398 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect -1916 549826 597980 549922
rect -1916 544350 597980 544446
rect -1916 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 3250 544350
rect 3306 544294 3374 544350
rect 3430 544294 3498 544350
rect 3554 544294 3622 544350
rect 3678 544294 21250 544350
rect 21306 544294 21374 544350
rect 21430 544294 21498 544350
rect 21554 544294 21622 544350
rect 21678 544294 39250 544350
rect 39306 544294 39374 544350
rect 39430 544294 39498 544350
rect 39554 544294 39622 544350
rect 39678 544294 57250 544350
rect 57306 544294 57374 544350
rect 57430 544294 57498 544350
rect 57554 544294 57622 544350
rect 57678 544294 75250 544350
rect 75306 544294 75374 544350
rect 75430 544294 75498 544350
rect 75554 544294 75622 544350
rect 75678 544294 93250 544350
rect 93306 544294 93374 544350
rect 93430 544294 93498 544350
rect 93554 544294 93622 544350
rect 93678 544294 111250 544350
rect 111306 544294 111374 544350
rect 111430 544294 111498 544350
rect 111554 544294 111622 544350
rect 111678 544294 129250 544350
rect 129306 544294 129374 544350
rect 129430 544294 129498 544350
rect 129554 544294 129622 544350
rect 129678 544294 147250 544350
rect 147306 544294 147374 544350
rect 147430 544294 147498 544350
rect 147554 544294 147622 544350
rect 147678 544294 165250 544350
rect 165306 544294 165374 544350
rect 165430 544294 165498 544350
rect 165554 544294 165622 544350
rect 165678 544294 183250 544350
rect 183306 544294 183374 544350
rect 183430 544294 183498 544350
rect 183554 544294 183622 544350
rect 183678 544294 201250 544350
rect 201306 544294 201374 544350
rect 201430 544294 201498 544350
rect 201554 544294 201622 544350
rect 201678 544294 219250 544350
rect 219306 544294 219374 544350
rect 219430 544294 219498 544350
rect 219554 544294 219622 544350
rect 219678 544294 237250 544350
rect 237306 544294 237374 544350
rect 237430 544294 237498 544350
rect 237554 544294 237622 544350
rect 237678 544294 255250 544350
rect 255306 544294 255374 544350
rect 255430 544294 255498 544350
rect 255554 544294 255622 544350
rect 255678 544294 273250 544350
rect 273306 544294 273374 544350
rect 273430 544294 273498 544350
rect 273554 544294 273622 544350
rect 273678 544294 291250 544350
rect 291306 544294 291374 544350
rect 291430 544294 291498 544350
rect 291554 544294 291622 544350
rect 291678 544294 309250 544350
rect 309306 544294 309374 544350
rect 309430 544294 309498 544350
rect 309554 544294 309622 544350
rect 309678 544294 327250 544350
rect 327306 544294 327374 544350
rect 327430 544294 327498 544350
rect 327554 544294 327622 544350
rect 327678 544294 345250 544350
rect 345306 544294 345374 544350
rect 345430 544294 345498 544350
rect 345554 544294 345622 544350
rect 345678 544294 363250 544350
rect 363306 544294 363374 544350
rect 363430 544294 363498 544350
rect 363554 544294 363622 544350
rect 363678 544294 381250 544350
rect 381306 544294 381374 544350
rect 381430 544294 381498 544350
rect 381554 544294 381622 544350
rect 381678 544294 399250 544350
rect 399306 544294 399374 544350
rect 399430 544294 399498 544350
rect 399554 544294 399622 544350
rect 399678 544294 417250 544350
rect 417306 544294 417374 544350
rect 417430 544294 417498 544350
rect 417554 544294 417622 544350
rect 417678 544294 435250 544350
rect 435306 544294 435374 544350
rect 435430 544294 435498 544350
rect 435554 544294 435622 544350
rect 435678 544294 453250 544350
rect 453306 544294 453374 544350
rect 453430 544294 453498 544350
rect 453554 544294 453622 544350
rect 453678 544294 471250 544350
rect 471306 544294 471374 544350
rect 471430 544294 471498 544350
rect 471554 544294 471622 544350
rect 471678 544294 489250 544350
rect 489306 544294 489374 544350
rect 489430 544294 489498 544350
rect 489554 544294 489622 544350
rect 489678 544294 507250 544350
rect 507306 544294 507374 544350
rect 507430 544294 507498 544350
rect 507554 544294 507622 544350
rect 507678 544294 525250 544350
rect 525306 544294 525374 544350
rect 525430 544294 525498 544350
rect 525554 544294 525622 544350
rect 525678 544294 543250 544350
rect 543306 544294 543374 544350
rect 543430 544294 543498 544350
rect 543554 544294 543622 544350
rect 543678 544294 561250 544350
rect 561306 544294 561374 544350
rect 561430 544294 561498 544350
rect 561554 544294 561622 544350
rect 561678 544294 579250 544350
rect 579306 544294 579374 544350
rect 579430 544294 579498 544350
rect 579554 544294 579622 544350
rect 579678 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597980 544350
rect -1916 544226 597980 544294
rect -1916 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 3250 544226
rect 3306 544170 3374 544226
rect 3430 544170 3498 544226
rect 3554 544170 3622 544226
rect 3678 544170 21250 544226
rect 21306 544170 21374 544226
rect 21430 544170 21498 544226
rect 21554 544170 21622 544226
rect 21678 544170 39250 544226
rect 39306 544170 39374 544226
rect 39430 544170 39498 544226
rect 39554 544170 39622 544226
rect 39678 544170 57250 544226
rect 57306 544170 57374 544226
rect 57430 544170 57498 544226
rect 57554 544170 57622 544226
rect 57678 544170 75250 544226
rect 75306 544170 75374 544226
rect 75430 544170 75498 544226
rect 75554 544170 75622 544226
rect 75678 544170 93250 544226
rect 93306 544170 93374 544226
rect 93430 544170 93498 544226
rect 93554 544170 93622 544226
rect 93678 544170 111250 544226
rect 111306 544170 111374 544226
rect 111430 544170 111498 544226
rect 111554 544170 111622 544226
rect 111678 544170 129250 544226
rect 129306 544170 129374 544226
rect 129430 544170 129498 544226
rect 129554 544170 129622 544226
rect 129678 544170 147250 544226
rect 147306 544170 147374 544226
rect 147430 544170 147498 544226
rect 147554 544170 147622 544226
rect 147678 544170 165250 544226
rect 165306 544170 165374 544226
rect 165430 544170 165498 544226
rect 165554 544170 165622 544226
rect 165678 544170 183250 544226
rect 183306 544170 183374 544226
rect 183430 544170 183498 544226
rect 183554 544170 183622 544226
rect 183678 544170 201250 544226
rect 201306 544170 201374 544226
rect 201430 544170 201498 544226
rect 201554 544170 201622 544226
rect 201678 544170 219250 544226
rect 219306 544170 219374 544226
rect 219430 544170 219498 544226
rect 219554 544170 219622 544226
rect 219678 544170 237250 544226
rect 237306 544170 237374 544226
rect 237430 544170 237498 544226
rect 237554 544170 237622 544226
rect 237678 544170 255250 544226
rect 255306 544170 255374 544226
rect 255430 544170 255498 544226
rect 255554 544170 255622 544226
rect 255678 544170 273250 544226
rect 273306 544170 273374 544226
rect 273430 544170 273498 544226
rect 273554 544170 273622 544226
rect 273678 544170 291250 544226
rect 291306 544170 291374 544226
rect 291430 544170 291498 544226
rect 291554 544170 291622 544226
rect 291678 544170 309250 544226
rect 309306 544170 309374 544226
rect 309430 544170 309498 544226
rect 309554 544170 309622 544226
rect 309678 544170 327250 544226
rect 327306 544170 327374 544226
rect 327430 544170 327498 544226
rect 327554 544170 327622 544226
rect 327678 544170 345250 544226
rect 345306 544170 345374 544226
rect 345430 544170 345498 544226
rect 345554 544170 345622 544226
rect 345678 544170 363250 544226
rect 363306 544170 363374 544226
rect 363430 544170 363498 544226
rect 363554 544170 363622 544226
rect 363678 544170 381250 544226
rect 381306 544170 381374 544226
rect 381430 544170 381498 544226
rect 381554 544170 381622 544226
rect 381678 544170 399250 544226
rect 399306 544170 399374 544226
rect 399430 544170 399498 544226
rect 399554 544170 399622 544226
rect 399678 544170 417250 544226
rect 417306 544170 417374 544226
rect 417430 544170 417498 544226
rect 417554 544170 417622 544226
rect 417678 544170 435250 544226
rect 435306 544170 435374 544226
rect 435430 544170 435498 544226
rect 435554 544170 435622 544226
rect 435678 544170 453250 544226
rect 453306 544170 453374 544226
rect 453430 544170 453498 544226
rect 453554 544170 453622 544226
rect 453678 544170 471250 544226
rect 471306 544170 471374 544226
rect 471430 544170 471498 544226
rect 471554 544170 471622 544226
rect 471678 544170 489250 544226
rect 489306 544170 489374 544226
rect 489430 544170 489498 544226
rect 489554 544170 489622 544226
rect 489678 544170 507250 544226
rect 507306 544170 507374 544226
rect 507430 544170 507498 544226
rect 507554 544170 507622 544226
rect 507678 544170 525250 544226
rect 525306 544170 525374 544226
rect 525430 544170 525498 544226
rect 525554 544170 525622 544226
rect 525678 544170 543250 544226
rect 543306 544170 543374 544226
rect 543430 544170 543498 544226
rect 543554 544170 543622 544226
rect 543678 544170 561250 544226
rect 561306 544170 561374 544226
rect 561430 544170 561498 544226
rect 561554 544170 561622 544226
rect 561678 544170 579250 544226
rect 579306 544170 579374 544226
rect 579430 544170 579498 544226
rect 579554 544170 579622 544226
rect 579678 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597980 544226
rect -1916 544102 597980 544170
rect -1916 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 3250 544102
rect 3306 544046 3374 544102
rect 3430 544046 3498 544102
rect 3554 544046 3622 544102
rect 3678 544046 21250 544102
rect 21306 544046 21374 544102
rect 21430 544046 21498 544102
rect 21554 544046 21622 544102
rect 21678 544046 39250 544102
rect 39306 544046 39374 544102
rect 39430 544046 39498 544102
rect 39554 544046 39622 544102
rect 39678 544046 57250 544102
rect 57306 544046 57374 544102
rect 57430 544046 57498 544102
rect 57554 544046 57622 544102
rect 57678 544046 75250 544102
rect 75306 544046 75374 544102
rect 75430 544046 75498 544102
rect 75554 544046 75622 544102
rect 75678 544046 93250 544102
rect 93306 544046 93374 544102
rect 93430 544046 93498 544102
rect 93554 544046 93622 544102
rect 93678 544046 111250 544102
rect 111306 544046 111374 544102
rect 111430 544046 111498 544102
rect 111554 544046 111622 544102
rect 111678 544046 129250 544102
rect 129306 544046 129374 544102
rect 129430 544046 129498 544102
rect 129554 544046 129622 544102
rect 129678 544046 147250 544102
rect 147306 544046 147374 544102
rect 147430 544046 147498 544102
rect 147554 544046 147622 544102
rect 147678 544046 165250 544102
rect 165306 544046 165374 544102
rect 165430 544046 165498 544102
rect 165554 544046 165622 544102
rect 165678 544046 183250 544102
rect 183306 544046 183374 544102
rect 183430 544046 183498 544102
rect 183554 544046 183622 544102
rect 183678 544046 201250 544102
rect 201306 544046 201374 544102
rect 201430 544046 201498 544102
rect 201554 544046 201622 544102
rect 201678 544046 219250 544102
rect 219306 544046 219374 544102
rect 219430 544046 219498 544102
rect 219554 544046 219622 544102
rect 219678 544046 237250 544102
rect 237306 544046 237374 544102
rect 237430 544046 237498 544102
rect 237554 544046 237622 544102
rect 237678 544046 255250 544102
rect 255306 544046 255374 544102
rect 255430 544046 255498 544102
rect 255554 544046 255622 544102
rect 255678 544046 273250 544102
rect 273306 544046 273374 544102
rect 273430 544046 273498 544102
rect 273554 544046 273622 544102
rect 273678 544046 291250 544102
rect 291306 544046 291374 544102
rect 291430 544046 291498 544102
rect 291554 544046 291622 544102
rect 291678 544046 309250 544102
rect 309306 544046 309374 544102
rect 309430 544046 309498 544102
rect 309554 544046 309622 544102
rect 309678 544046 327250 544102
rect 327306 544046 327374 544102
rect 327430 544046 327498 544102
rect 327554 544046 327622 544102
rect 327678 544046 345250 544102
rect 345306 544046 345374 544102
rect 345430 544046 345498 544102
rect 345554 544046 345622 544102
rect 345678 544046 363250 544102
rect 363306 544046 363374 544102
rect 363430 544046 363498 544102
rect 363554 544046 363622 544102
rect 363678 544046 381250 544102
rect 381306 544046 381374 544102
rect 381430 544046 381498 544102
rect 381554 544046 381622 544102
rect 381678 544046 399250 544102
rect 399306 544046 399374 544102
rect 399430 544046 399498 544102
rect 399554 544046 399622 544102
rect 399678 544046 417250 544102
rect 417306 544046 417374 544102
rect 417430 544046 417498 544102
rect 417554 544046 417622 544102
rect 417678 544046 435250 544102
rect 435306 544046 435374 544102
rect 435430 544046 435498 544102
rect 435554 544046 435622 544102
rect 435678 544046 453250 544102
rect 453306 544046 453374 544102
rect 453430 544046 453498 544102
rect 453554 544046 453622 544102
rect 453678 544046 471250 544102
rect 471306 544046 471374 544102
rect 471430 544046 471498 544102
rect 471554 544046 471622 544102
rect 471678 544046 489250 544102
rect 489306 544046 489374 544102
rect 489430 544046 489498 544102
rect 489554 544046 489622 544102
rect 489678 544046 507250 544102
rect 507306 544046 507374 544102
rect 507430 544046 507498 544102
rect 507554 544046 507622 544102
rect 507678 544046 525250 544102
rect 525306 544046 525374 544102
rect 525430 544046 525498 544102
rect 525554 544046 525622 544102
rect 525678 544046 543250 544102
rect 543306 544046 543374 544102
rect 543430 544046 543498 544102
rect 543554 544046 543622 544102
rect 543678 544046 561250 544102
rect 561306 544046 561374 544102
rect 561430 544046 561498 544102
rect 561554 544046 561622 544102
rect 561678 544046 579250 544102
rect 579306 544046 579374 544102
rect 579430 544046 579498 544102
rect 579554 544046 579622 544102
rect 579678 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597980 544102
rect -1916 543978 597980 544046
rect -1916 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 3250 543978
rect 3306 543922 3374 543978
rect 3430 543922 3498 543978
rect 3554 543922 3622 543978
rect 3678 543922 21250 543978
rect 21306 543922 21374 543978
rect 21430 543922 21498 543978
rect 21554 543922 21622 543978
rect 21678 543922 39250 543978
rect 39306 543922 39374 543978
rect 39430 543922 39498 543978
rect 39554 543922 39622 543978
rect 39678 543922 57250 543978
rect 57306 543922 57374 543978
rect 57430 543922 57498 543978
rect 57554 543922 57622 543978
rect 57678 543922 75250 543978
rect 75306 543922 75374 543978
rect 75430 543922 75498 543978
rect 75554 543922 75622 543978
rect 75678 543922 93250 543978
rect 93306 543922 93374 543978
rect 93430 543922 93498 543978
rect 93554 543922 93622 543978
rect 93678 543922 111250 543978
rect 111306 543922 111374 543978
rect 111430 543922 111498 543978
rect 111554 543922 111622 543978
rect 111678 543922 129250 543978
rect 129306 543922 129374 543978
rect 129430 543922 129498 543978
rect 129554 543922 129622 543978
rect 129678 543922 147250 543978
rect 147306 543922 147374 543978
rect 147430 543922 147498 543978
rect 147554 543922 147622 543978
rect 147678 543922 165250 543978
rect 165306 543922 165374 543978
rect 165430 543922 165498 543978
rect 165554 543922 165622 543978
rect 165678 543922 183250 543978
rect 183306 543922 183374 543978
rect 183430 543922 183498 543978
rect 183554 543922 183622 543978
rect 183678 543922 201250 543978
rect 201306 543922 201374 543978
rect 201430 543922 201498 543978
rect 201554 543922 201622 543978
rect 201678 543922 219250 543978
rect 219306 543922 219374 543978
rect 219430 543922 219498 543978
rect 219554 543922 219622 543978
rect 219678 543922 237250 543978
rect 237306 543922 237374 543978
rect 237430 543922 237498 543978
rect 237554 543922 237622 543978
rect 237678 543922 255250 543978
rect 255306 543922 255374 543978
rect 255430 543922 255498 543978
rect 255554 543922 255622 543978
rect 255678 543922 273250 543978
rect 273306 543922 273374 543978
rect 273430 543922 273498 543978
rect 273554 543922 273622 543978
rect 273678 543922 291250 543978
rect 291306 543922 291374 543978
rect 291430 543922 291498 543978
rect 291554 543922 291622 543978
rect 291678 543922 309250 543978
rect 309306 543922 309374 543978
rect 309430 543922 309498 543978
rect 309554 543922 309622 543978
rect 309678 543922 327250 543978
rect 327306 543922 327374 543978
rect 327430 543922 327498 543978
rect 327554 543922 327622 543978
rect 327678 543922 345250 543978
rect 345306 543922 345374 543978
rect 345430 543922 345498 543978
rect 345554 543922 345622 543978
rect 345678 543922 363250 543978
rect 363306 543922 363374 543978
rect 363430 543922 363498 543978
rect 363554 543922 363622 543978
rect 363678 543922 381250 543978
rect 381306 543922 381374 543978
rect 381430 543922 381498 543978
rect 381554 543922 381622 543978
rect 381678 543922 399250 543978
rect 399306 543922 399374 543978
rect 399430 543922 399498 543978
rect 399554 543922 399622 543978
rect 399678 543922 417250 543978
rect 417306 543922 417374 543978
rect 417430 543922 417498 543978
rect 417554 543922 417622 543978
rect 417678 543922 435250 543978
rect 435306 543922 435374 543978
rect 435430 543922 435498 543978
rect 435554 543922 435622 543978
rect 435678 543922 453250 543978
rect 453306 543922 453374 543978
rect 453430 543922 453498 543978
rect 453554 543922 453622 543978
rect 453678 543922 471250 543978
rect 471306 543922 471374 543978
rect 471430 543922 471498 543978
rect 471554 543922 471622 543978
rect 471678 543922 489250 543978
rect 489306 543922 489374 543978
rect 489430 543922 489498 543978
rect 489554 543922 489622 543978
rect 489678 543922 507250 543978
rect 507306 543922 507374 543978
rect 507430 543922 507498 543978
rect 507554 543922 507622 543978
rect 507678 543922 525250 543978
rect 525306 543922 525374 543978
rect 525430 543922 525498 543978
rect 525554 543922 525622 543978
rect 525678 543922 543250 543978
rect 543306 543922 543374 543978
rect 543430 543922 543498 543978
rect 543554 543922 543622 543978
rect 543678 543922 561250 543978
rect 561306 543922 561374 543978
rect 561430 543922 561498 543978
rect 561554 543922 561622 543978
rect 561678 543922 579250 543978
rect 579306 543922 579374 543978
rect 579430 543922 579498 543978
rect 579554 543922 579622 543978
rect 579678 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597980 543978
rect -1916 543826 597980 543922
rect -1916 532350 597980 532446
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 6970 532350
rect 7026 532294 7094 532350
rect 7150 532294 7218 532350
rect 7274 532294 7342 532350
rect 7398 532294 24970 532350
rect 25026 532294 25094 532350
rect 25150 532294 25218 532350
rect 25274 532294 25342 532350
rect 25398 532294 42970 532350
rect 43026 532294 43094 532350
rect 43150 532294 43218 532350
rect 43274 532294 43342 532350
rect 43398 532294 60970 532350
rect 61026 532294 61094 532350
rect 61150 532294 61218 532350
rect 61274 532294 61342 532350
rect 61398 532294 78970 532350
rect 79026 532294 79094 532350
rect 79150 532294 79218 532350
rect 79274 532294 79342 532350
rect 79398 532294 96970 532350
rect 97026 532294 97094 532350
rect 97150 532294 97218 532350
rect 97274 532294 97342 532350
rect 97398 532294 114970 532350
rect 115026 532294 115094 532350
rect 115150 532294 115218 532350
rect 115274 532294 115342 532350
rect 115398 532294 132970 532350
rect 133026 532294 133094 532350
rect 133150 532294 133218 532350
rect 133274 532294 133342 532350
rect 133398 532294 150970 532350
rect 151026 532294 151094 532350
rect 151150 532294 151218 532350
rect 151274 532294 151342 532350
rect 151398 532294 168970 532350
rect 169026 532294 169094 532350
rect 169150 532294 169218 532350
rect 169274 532294 169342 532350
rect 169398 532294 186970 532350
rect 187026 532294 187094 532350
rect 187150 532294 187218 532350
rect 187274 532294 187342 532350
rect 187398 532294 204970 532350
rect 205026 532294 205094 532350
rect 205150 532294 205218 532350
rect 205274 532294 205342 532350
rect 205398 532294 222970 532350
rect 223026 532294 223094 532350
rect 223150 532294 223218 532350
rect 223274 532294 223342 532350
rect 223398 532294 240970 532350
rect 241026 532294 241094 532350
rect 241150 532294 241218 532350
rect 241274 532294 241342 532350
rect 241398 532294 258970 532350
rect 259026 532294 259094 532350
rect 259150 532294 259218 532350
rect 259274 532294 259342 532350
rect 259398 532294 276970 532350
rect 277026 532294 277094 532350
rect 277150 532294 277218 532350
rect 277274 532294 277342 532350
rect 277398 532294 294970 532350
rect 295026 532294 295094 532350
rect 295150 532294 295218 532350
rect 295274 532294 295342 532350
rect 295398 532294 312970 532350
rect 313026 532294 313094 532350
rect 313150 532294 313218 532350
rect 313274 532294 313342 532350
rect 313398 532294 330970 532350
rect 331026 532294 331094 532350
rect 331150 532294 331218 532350
rect 331274 532294 331342 532350
rect 331398 532294 348970 532350
rect 349026 532294 349094 532350
rect 349150 532294 349218 532350
rect 349274 532294 349342 532350
rect 349398 532294 366970 532350
rect 367026 532294 367094 532350
rect 367150 532294 367218 532350
rect 367274 532294 367342 532350
rect 367398 532294 384970 532350
rect 385026 532294 385094 532350
rect 385150 532294 385218 532350
rect 385274 532294 385342 532350
rect 385398 532294 402970 532350
rect 403026 532294 403094 532350
rect 403150 532294 403218 532350
rect 403274 532294 403342 532350
rect 403398 532294 420970 532350
rect 421026 532294 421094 532350
rect 421150 532294 421218 532350
rect 421274 532294 421342 532350
rect 421398 532294 438970 532350
rect 439026 532294 439094 532350
rect 439150 532294 439218 532350
rect 439274 532294 439342 532350
rect 439398 532294 456970 532350
rect 457026 532294 457094 532350
rect 457150 532294 457218 532350
rect 457274 532294 457342 532350
rect 457398 532294 474970 532350
rect 475026 532294 475094 532350
rect 475150 532294 475218 532350
rect 475274 532294 475342 532350
rect 475398 532294 492970 532350
rect 493026 532294 493094 532350
rect 493150 532294 493218 532350
rect 493274 532294 493342 532350
rect 493398 532294 510970 532350
rect 511026 532294 511094 532350
rect 511150 532294 511218 532350
rect 511274 532294 511342 532350
rect 511398 532294 528970 532350
rect 529026 532294 529094 532350
rect 529150 532294 529218 532350
rect 529274 532294 529342 532350
rect 529398 532294 546970 532350
rect 547026 532294 547094 532350
rect 547150 532294 547218 532350
rect 547274 532294 547342 532350
rect 547398 532294 564970 532350
rect 565026 532294 565094 532350
rect 565150 532294 565218 532350
rect 565274 532294 565342 532350
rect 565398 532294 582970 532350
rect 583026 532294 583094 532350
rect 583150 532294 583218 532350
rect 583274 532294 583342 532350
rect 583398 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect -1916 532226 597980 532294
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 6970 532226
rect 7026 532170 7094 532226
rect 7150 532170 7218 532226
rect 7274 532170 7342 532226
rect 7398 532170 24970 532226
rect 25026 532170 25094 532226
rect 25150 532170 25218 532226
rect 25274 532170 25342 532226
rect 25398 532170 42970 532226
rect 43026 532170 43094 532226
rect 43150 532170 43218 532226
rect 43274 532170 43342 532226
rect 43398 532170 60970 532226
rect 61026 532170 61094 532226
rect 61150 532170 61218 532226
rect 61274 532170 61342 532226
rect 61398 532170 78970 532226
rect 79026 532170 79094 532226
rect 79150 532170 79218 532226
rect 79274 532170 79342 532226
rect 79398 532170 96970 532226
rect 97026 532170 97094 532226
rect 97150 532170 97218 532226
rect 97274 532170 97342 532226
rect 97398 532170 114970 532226
rect 115026 532170 115094 532226
rect 115150 532170 115218 532226
rect 115274 532170 115342 532226
rect 115398 532170 132970 532226
rect 133026 532170 133094 532226
rect 133150 532170 133218 532226
rect 133274 532170 133342 532226
rect 133398 532170 150970 532226
rect 151026 532170 151094 532226
rect 151150 532170 151218 532226
rect 151274 532170 151342 532226
rect 151398 532170 168970 532226
rect 169026 532170 169094 532226
rect 169150 532170 169218 532226
rect 169274 532170 169342 532226
rect 169398 532170 186970 532226
rect 187026 532170 187094 532226
rect 187150 532170 187218 532226
rect 187274 532170 187342 532226
rect 187398 532170 204970 532226
rect 205026 532170 205094 532226
rect 205150 532170 205218 532226
rect 205274 532170 205342 532226
rect 205398 532170 222970 532226
rect 223026 532170 223094 532226
rect 223150 532170 223218 532226
rect 223274 532170 223342 532226
rect 223398 532170 240970 532226
rect 241026 532170 241094 532226
rect 241150 532170 241218 532226
rect 241274 532170 241342 532226
rect 241398 532170 258970 532226
rect 259026 532170 259094 532226
rect 259150 532170 259218 532226
rect 259274 532170 259342 532226
rect 259398 532170 276970 532226
rect 277026 532170 277094 532226
rect 277150 532170 277218 532226
rect 277274 532170 277342 532226
rect 277398 532170 294970 532226
rect 295026 532170 295094 532226
rect 295150 532170 295218 532226
rect 295274 532170 295342 532226
rect 295398 532170 312970 532226
rect 313026 532170 313094 532226
rect 313150 532170 313218 532226
rect 313274 532170 313342 532226
rect 313398 532170 330970 532226
rect 331026 532170 331094 532226
rect 331150 532170 331218 532226
rect 331274 532170 331342 532226
rect 331398 532170 348970 532226
rect 349026 532170 349094 532226
rect 349150 532170 349218 532226
rect 349274 532170 349342 532226
rect 349398 532170 366970 532226
rect 367026 532170 367094 532226
rect 367150 532170 367218 532226
rect 367274 532170 367342 532226
rect 367398 532170 384970 532226
rect 385026 532170 385094 532226
rect 385150 532170 385218 532226
rect 385274 532170 385342 532226
rect 385398 532170 402970 532226
rect 403026 532170 403094 532226
rect 403150 532170 403218 532226
rect 403274 532170 403342 532226
rect 403398 532170 420970 532226
rect 421026 532170 421094 532226
rect 421150 532170 421218 532226
rect 421274 532170 421342 532226
rect 421398 532170 438970 532226
rect 439026 532170 439094 532226
rect 439150 532170 439218 532226
rect 439274 532170 439342 532226
rect 439398 532170 456970 532226
rect 457026 532170 457094 532226
rect 457150 532170 457218 532226
rect 457274 532170 457342 532226
rect 457398 532170 474970 532226
rect 475026 532170 475094 532226
rect 475150 532170 475218 532226
rect 475274 532170 475342 532226
rect 475398 532170 492970 532226
rect 493026 532170 493094 532226
rect 493150 532170 493218 532226
rect 493274 532170 493342 532226
rect 493398 532170 510970 532226
rect 511026 532170 511094 532226
rect 511150 532170 511218 532226
rect 511274 532170 511342 532226
rect 511398 532170 528970 532226
rect 529026 532170 529094 532226
rect 529150 532170 529218 532226
rect 529274 532170 529342 532226
rect 529398 532170 546970 532226
rect 547026 532170 547094 532226
rect 547150 532170 547218 532226
rect 547274 532170 547342 532226
rect 547398 532170 564970 532226
rect 565026 532170 565094 532226
rect 565150 532170 565218 532226
rect 565274 532170 565342 532226
rect 565398 532170 582970 532226
rect 583026 532170 583094 532226
rect 583150 532170 583218 532226
rect 583274 532170 583342 532226
rect 583398 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect -1916 532102 597980 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 6970 532102
rect 7026 532046 7094 532102
rect 7150 532046 7218 532102
rect 7274 532046 7342 532102
rect 7398 532046 24970 532102
rect 25026 532046 25094 532102
rect 25150 532046 25218 532102
rect 25274 532046 25342 532102
rect 25398 532046 42970 532102
rect 43026 532046 43094 532102
rect 43150 532046 43218 532102
rect 43274 532046 43342 532102
rect 43398 532046 60970 532102
rect 61026 532046 61094 532102
rect 61150 532046 61218 532102
rect 61274 532046 61342 532102
rect 61398 532046 78970 532102
rect 79026 532046 79094 532102
rect 79150 532046 79218 532102
rect 79274 532046 79342 532102
rect 79398 532046 96970 532102
rect 97026 532046 97094 532102
rect 97150 532046 97218 532102
rect 97274 532046 97342 532102
rect 97398 532046 114970 532102
rect 115026 532046 115094 532102
rect 115150 532046 115218 532102
rect 115274 532046 115342 532102
rect 115398 532046 132970 532102
rect 133026 532046 133094 532102
rect 133150 532046 133218 532102
rect 133274 532046 133342 532102
rect 133398 532046 150970 532102
rect 151026 532046 151094 532102
rect 151150 532046 151218 532102
rect 151274 532046 151342 532102
rect 151398 532046 168970 532102
rect 169026 532046 169094 532102
rect 169150 532046 169218 532102
rect 169274 532046 169342 532102
rect 169398 532046 186970 532102
rect 187026 532046 187094 532102
rect 187150 532046 187218 532102
rect 187274 532046 187342 532102
rect 187398 532046 204970 532102
rect 205026 532046 205094 532102
rect 205150 532046 205218 532102
rect 205274 532046 205342 532102
rect 205398 532046 222970 532102
rect 223026 532046 223094 532102
rect 223150 532046 223218 532102
rect 223274 532046 223342 532102
rect 223398 532046 240970 532102
rect 241026 532046 241094 532102
rect 241150 532046 241218 532102
rect 241274 532046 241342 532102
rect 241398 532046 258970 532102
rect 259026 532046 259094 532102
rect 259150 532046 259218 532102
rect 259274 532046 259342 532102
rect 259398 532046 276970 532102
rect 277026 532046 277094 532102
rect 277150 532046 277218 532102
rect 277274 532046 277342 532102
rect 277398 532046 294970 532102
rect 295026 532046 295094 532102
rect 295150 532046 295218 532102
rect 295274 532046 295342 532102
rect 295398 532046 312970 532102
rect 313026 532046 313094 532102
rect 313150 532046 313218 532102
rect 313274 532046 313342 532102
rect 313398 532046 330970 532102
rect 331026 532046 331094 532102
rect 331150 532046 331218 532102
rect 331274 532046 331342 532102
rect 331398 532046 348970 532102
rect 349026 532046 349094 532102
rect 349150 532046 349218 532102
rect 349274 532046 349342 532102
rect 349398 532046 366970 532102
rect 367026 532046 367094 532102
rect 367150 532046 367218 532102
rect 367274 532046 367342 532102
rect 367398 532046 384970 532102
rect 385026 532046 385094 532102
rect 385150 532046 385218 532102
rect 385274 532046 385342 532102
rect 385398 532046 402970 532102
rect 403026 532046 403094 532102
rect 403150 532046 403218 532102
rect 403274 532046 403342 532102
rect 403398 532046 420970 532102
rect 421026 532046 421094 532102
rect 421150 532046 421218 532102
rect 421274 532046 421342 532102
rect 421398 532046 438970 532102
rect 439026 532046 439094 532102
rect 439150 532046 439218 532102
rect 439274 532046 439342 532102
rect 439398 532046 456970 532102
rect 457026 532046 457094 532102
rect 457150 532046 457218 532102
rect 457274 532046 457342 532102
rect 457398 532046 474970 532102
rect 475026 532046 475094 532102
rect 475150 532046 475218 532102
rect 475274 532046 475342 532102
rect 475398 532046 492970 532102
rect 493026 532046 493094 532102
rect 493150 532046 493218 532102
rect 493274 532046 493342 532102
rect 493398 532046 510970 532102
rect 511026 532046 511094 532102
rect 511150 532046 511218 532102
rect 511274 532046 511342 532102
rect 511398 532046 528970 532102
rect 529026 532046 529094 532102
rect 529150 532046 529218 532102
rect 529274 532046 529342 532102
rect 529398 532046 546970 532102
rect 547026 532046 547094 532102
rect 547150 532046 547218 532102
rect 547274 532046 547342 532102
rect 547398 532046 564970 532102
rect 565026 532046 565094 532102
rect 565150 532046 565218 532102
rect 565274 532046 565342 532102
rect 565398 532046 582970 532102
rect 583026 532046 583094 532102
rect 583150 532046 583218 532102
rect 583274 532046 583342 532102
rect 583398 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect -1916 531978 597980 532046
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 6970 531978
rect 7026 531922 7094 531978
rect 7150 531922 7218 531978
rect 7274 531922 7342 531978
rect 7398 531922 24970 531978
rect 25026 531922 25094 531978
rect 25150 531922 25218 531978
rect 25274 531922 25342 531978
rect 25398 531922 42970 531978
rect 43026 531922 43094 531978
rect 43150 531922 43218 531978
rect 43274 531922 43342 531978
rect 43398 531922 60970 531978
rect 61026 531922 61094 531978
rect 61150 531922 61218 531978
rect 61274 531922 61342 531978
rect 61398 531922 78970 531978
rect 79026 531922 79094 531978
rect 79150 531922 79218 531978
rect 79274 531922 79342 531978
rect 79398 531922 96970 531978
rect 97026 531922 97094 531978
rect 97150 531922 97218 531978
rect 97274 531922 97342 531978
rect 97398 531922 114970 531978
rect 115026 531922 115094 531978
rect 115150 531922 115218 531978
rect 115274 531922 115342 531978
rect 115398 531922 132970 531978
rect 133026 531922 133094 531978
rect 133150 531922 133218 531978
rect 133274 531922 133342 531978
rect 133398 531922 150970 531978
rect 151026 531922 151094 531978
rect 151150 531922 151218 531978
rect 151274 531922 151342 531978
rect 151398 531922 168970 531978
rect 169026 531922 169094 531978
rect 169150 531922 169218 531978
rect 169274 531922 169342 531978
rect 169398 531922 186970 531978
rect 187026 531922 187094 531978
rect 187150 531922 187218 531978
rect 187274 531922 187342 531978
rect 187398 531922 204970 531978
rect 205026 531922 205094 531978
rect 205150 531922 205218 531978
rect 205274 531922 205342 531978
rect 205398 531922 222970 531978
rect 223026 531922 223094 531978
rect 223150 531922 223218 531978
rect 223274 531922 223342 531978
rect 223398 531922 240970 531978
rect 241026 531922 241094 531978
rect 241150 531922 241218 531978
rect 241274 531922 241342 531978
rect 241398 531922 258970 531978
rect 259026 531922 259094 531978
rect 259150 531922 259218 531978
rect 259274 531922 259342 531978
rect 259398 531922 276970 531978
rect 277026 531922 277094 531978
rect 277150 531922 277218 531978
rect 277274 531922 277342 531978
rect 277398 531922 294970 531978
rect 295026 531922 295094 531978
rect 295150 531922 295218 531978
rect 295274 531922 295342 531978
rect 295398 531922 312970 531978
rect 313026 531922 313094 531978
rect 313150 531922 313218 531978
rect 313274 531922 313342 531978
rect 313398 531922 330970 531978
rect 331026 531922 331094 531978
rect 331150 531922 331218 531978
rect 331274 531922 331342 531978
rect 331398 531922 348970 531978
rect 349026 531922 349094 531978
rect 349150 531922 349218 531978
rect 349274 531922 349342 531978
rect 349398 531922 366970 531978
rect 367026 531922 367094 531978
rect 367150 531922 367218 531978
rect 367274 531922 367342 531978
rect 367398 531922 384970 531978
rect 385026 531922 385094 531978
rect 385150 531922 385218 531978
rect 385274 531922 385342 531978
rect 385398 531922 402970 531978
rect 403026 531922 403094 531978
rect 403150 531922 403218 531978
rect 403274 531922 403342 531978
rect 403398 531922 420970 531978
rect 421026 531922 421094 531978
rect 421150 531922 421218 531978
rect 421274 531922 421342 531978
rect 421398 531922 438970 531978
rect 439026 531922 439094 531978
rect 439150 531922 439218 531978
rect 439274 531922 439342 531978
rect 439398 531922 456970 531978
rect 457026 531922 457094 531978
rect 457150 531922 457218 531978
rect 457274 531922 457342 531978
rect 457398 531922 474970 531978
rect 475026 531922 475094 531978
rect 475150 531922 475218 531978
rect 475274 531922 475342 531978
rect 475398 531922 492970 531978
rect 493026 531922 493094 531978
rect 493150 531922 493218 531978
rect 493274 531922 493342 531978
rect 493398 531922 510970 531978
rect 511026 531922 511094 531978
rect 511150 531922 511218 531978
rect 511274 531922 511342 531978
rect 511398 531922 528970 531978
rect 529026 531922 529094 531978
rect 529150 531922 529218 531978
rect 529274 531922 529342 531978
rect 529398 531922 546970 531978
rect 547026 531922 547094 531978
rect 547150 531922 547218 531978
rect 547274 531922 547342 531978
rect 547398 531922 564970 531978
rect 565026 531922 565094 531978
rect 565150 531922 565218 531978
rect 565274 531922 565342 531978
rect 565398 531922 582970 531978
rect 583026 531922 583094 531978
rect 583150 531922 583218 531978
rect 583274 531922 583342 531978
rect 583398 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect -1916 531826 597980 531922
rect -1916 526350 597980 526446
rect -1916 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 3250 526350
rect 3306 526294 3374 526350
rect 3430 526294 3498 526350
rect 3554 526294 3622 526350
rect 3678 526294 21250 526350
rect 21306 526294 21374 526350
rect 21430 526294 21498 526350
rect 21554 526294 21622 526350
rect 21678 526294 39250 526350
rect 39306 526294 39374 526350
rect 39430 526294 39498 526350
rect 39554 526294 39622 526350
rect 39678 526294 57250 526350
rect 57306 526294 57374 526350
rect 57430 526294 57498 526350
rect 57554 526294 57622 526350
rect 57678 526294 75250 526350
rect 75306 526294 75374 526350
rect 75430 526294 75498 526350
rect 75554 526294 75622 526350
rect 75678 526294 93250 526350
rect 93306 526294 93374 526350
rect 93430 526294 93498 526350
rect 93554 526294 93622 526350
rect 93678 526294 111250 526350
rect 111306 526294 111374 526350
rect 111430 526294 111498 526350
rect 111554 526294 111622 526350
rect 111678 526294 561250 526350
rect 561306 526294 561374 526350
rect 561430 526294 561498 526350
rect 561554 526294 561622 526350
rect 561678 526294 579250 526350
rect 579306 526294 579374 526350
rect 579430 526294 579498 526350
rect 579554 526294 579622 526350
rect 579678 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597980 526350
rect -1916 526293 597980 526294
rect -1916 526237 54518 526293
rect 54574 526237 54642 526293
rect 54698 526237 85238 526293
rect 85294 526237 85362 526293
rect 85418 526237 115958 526293
rect 116014 526237 116082 526293
rect 116138 526237 146678 526293
rect 146734 526237 146802 526293
rect 146858 526237 177398 526293
rect 177454 526237 177522 526293
rect 177578 526237 208118 526293
rect 208174 526237 208242 526293
rect 208298 526237 238838 526293
rect 238894 526237 238962 526293
rect 239018 526237 269558 526293
rect 269614 526237 269682 526293
rect 269738 526237 300278 526293
rect 300334 526237 300402 526293
rect 300458 526237 330998 526293
rect 331054 526237 331122 526293
rect 331178 526237 361718 526293
rect 361774 526237 361842 526293
rect 361898 526237 392438 526293
rect 392494 526237 392562 526293
rect 392618 526237 423158 526293
rect 423214 526237 423282 526293
rect 423338 526237 453878 526293
rect 453934 526237 454002 526293
rect 454058 526237 484598 526293
rect 484654 526237 484722 526293
rect 484778 526237 515318 526293
rect 515374 526237 515442 526293
rect 515498 526237 546038 526293
rect 546094 526237 546162 526293
rect 546218 526237 597980 526293
rect -1916 526226 597980 526237
rect -1916 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 3250 526226
rect 3306 526170 3374 526226
rect 3430 526170 3498 526226
rect 3554 526170 3622 526226
rect 3678 526170 21250 526226
rect 21306 526170 21374 526226
rect 21430 526170 21498 526226
rect 21554 526170 21622 526226
rect 21678 526170 39250 526226
rect 39306 526170 39374 526226
rect 39430 526170 39498 526226
rect 39554 526170 39622 526226
rect 39678 526170 57250 526226
rect 57306 526170 57374 526226
rect 57430 526170 57498 526226
rect 57554 526170 57622 526226
rect 57678 526170 75250 526226
rect 75306 526170 75374 526226
rect 75430 526170 75498 526226
rect 75554 526170 75622 526226
rect 75678 526170 93250 526226
rect 93306 526170 93374 526226
rect 93430 526170 93498 526226
rect 93554 526170 93622 526226
rect 93678 526170 111250 526226
rect 111306 526170 111374 526226
rect 111430 526170 111498 526226
rect 111554 526170 111622 526226
rect 111678 526170 561250 526226
rect 561306 526170 561374 526226
rect 561430 526170 561498 526226
rect 561554 526170 561622 526226
rect 561678 526170 579250 526226
rect 579306 526170 579374 526226
rect 579430 526170 579498 526226
rect 579554 526170 579622 526226
rect 579678 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597980 526226
rect -1916 526169 597980 526170
rect -1916 526113 54518 526169
rect 54574 526113 54642 526169
rect 54698 526113 85238 526169
rect 85294 526113 85362 526169
rect 85418 526113 115958 526169
rect 116014 526113 116082 526169
rect 116138 526113 146678 526169
rect 146734 526113 146802 526169
rect 146858 526113 177398 526169
rect 177454 526113 177522 526169
rect 177578 526113 208118 526169
rect 208174 526113 208242 526169
rect 208298 526113 238838 526169
rect 238894 526113 238962 526169
rect 239018 526113 269558 526169
rect 269614 526113 269682 526169
rect 269738 526113 300278 526169
rect 300334 526113 300402 526169
rect 300458 526113 330998 526169
rect 331054 526113 331122 526169
rect 331178 526113 361718 526169
rect 361774 526113 361842 526169
rect 361898 526113 392438 526169
rect 392494 526113 392562 526169
rect 392618 526113 423158 526169
rect 423214 526113 423282 526169
rect 423338 526113 453878 526169
rect 453934 526113 454002 526169
rect 454058 526113 484598 526169
rect 484654 526113 484722 526169
rect 484778 526113 515318 526169
rect 515374 526113 515442 526169
rect 515498 526113 546038 526169
rect 546094 526113 546162 526169
rect 546218 526113 597980 526169
rect -1916 526102 597980 526113
rect -1916 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 3250 526102
rect 3306 526046 3374 526102
rect 3430 526046 3498 526102
rect 3554 526046 3622 526102
rect 3678 526046 21250 526102
rect 21306 526046 21374 526102
rect 21430 526046 21498 526102
rect 21554 526046 21622 526102
rect 21678 526046 39250 526102
rect 39306 526046 39374 526102
rect 39430 526046 39498 526102
rect 39554 526046 39622 526102
rect 39678 526046 57250 526102
rect 57306 526046 57374 526102
rect 57430 526046 57498 526102
rect 57554 526046 57622 526102
rect 57678 526046 75250 526102
rect 75306 526046 75374 526102
rect 75430 526046 75498 526102
rect 75554 526046 75622 526102
rect 75678 526046 93250 526102
rect 93306 526046 93374 526102
rect 93430 526046 93498 526102
rect 93554 526046 93622 526102
rect 93678 526046 111250 526102
rect 111306 526046 111374 526102
rect 111430 526046 111498 526102
rect 111554 526046 111622 526102
rect 111678 526046 561250 526102
rect 561306 526046 561374 526102
rect 561430 526046 561498 526102
rect 561554 526046 561622 526102
rect 561678 526046 579250 526102
rect 579306 526046 579374 526102
rect 579430 526046 579498 526102
rect 579554 526046 579622 526102
rect 579678 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597980 526102
rect -1916 526045 597980 526046
rect -1916 525989 54518 526045
rect 54574 525989 54642 526045
rect 54698 525989 85238 526045
rect 85294 525989 85362 526045
rect 85418 525989 115958 526045
rect 116014 525989 116082 526045
rect 116138 525989 146678 526045
rect 146734 525989 146802 526045
rect 146858 525989 177398 526045
rect 177454 525989 177522 526045
rect 177578 525989 208118 526045
rect 208174 525989 208242 526045
rect 208298 525989 238838 526045
rect 238894 525989 238962 526045
rect 239018 525989 269558 526045
rect 269614 525989 269682 526045
rect 269738 525989 300278 526045
rect 300334 525989 300402 526045
rect 300458 525989 330998 526045
rect 331054 525989 331122 526045
rect 331178 525989 361718 526045
rect 361774 525989 361842 526045
rect 361898 525989 392438 526045
rect 392494 525989 392562 526045
rect 392618 525989 423158 526045
rect 423214 525989 423282 526045
rect 423338 525989 453878 526045
rect 453934 525989 454002 526045
rect 454058 525989 484598 526045
rect 484654 525989 484722 526045
rect 484778 525989 515318 526045
rect 515374 525989 515442 526045
rect 515498 525989 546038 526045
rect 546094 525989 546162 526045
rect 546218 525989 597980 526045
rect -1916 525978 597980 525989
rect -1916 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 3250 525978
rect 3306 525922 3374 525978
rect 3430 525922 3498 525978
rect 3554 525922 3622 525978
rect 3678 525922 21250 525978
rect 21306 525922 21374 525978
rect 21430 525922 21498 525978
rect 21554 525922 21622 525978
rect 21678 525922 39250 525978
rect 39306 525922 39374 525978
rect 39430 525922 39498 525978
rect 39554 525922 39622 525978
rect 39678 525922 57250 525978
rect 57306 525922 57374 525978
rect 57430 525922 57498 525978
rect 57554 525922 57622 525978
rect 57678 525922 75250 525978
rect 75306 525922 75374 525978
rect 75430 525922 75498 525978
rect 75554 525922 75622 525978
rect 75678 525922 93250 525978
rect 93306 525922 93374 525978
rect 93430 525922 93498 525978
rect 93554 525922 93622 525978
rect 93678 525922 111250 525978
rect 111306 525922 111374 525978
rect 111430 525922 111498 525978
rect 111554 525922 111622 525978
rect 111678 525922 561250 525978
rect 561306 525922 561374 525978
rect 561430 525922 561498 525978
rect 561554 525922 561622 525978
rect 561678 525922 579250 525978
rect 579306 525922 579374 525978
rect 579430 525922 579498 525978
rect 579554 525922 579622 525978
rect 579678 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597980 525978
rect -1916 525921 597980 525922
rect -1916 525865 54518 525921
rect 54574 525865 54642 525921
rect 54698 525865 85238 525921
rect 85294 525865 85362 525921
rect 85418 525865 115958 525921
rect 116014 525865 116082 525921
rect 116138 525865 146678 525921
rect 146734 525865 146802 525921
rect 146858 525865 177398 525921
rect 177454 525865 177522 525921
rect 177578 525865 208118 525921
rect 208174 525865 208242 525921
rect 208298 525865 238838 525921
rect 238894 525865 238962 525921
rect 239018 525865 269558 525921
rect 269614 525865 269682 525921
rect 269738 525865 300278 525921
rect 300334 525865 300402 525921
rect 300458 525865 330998 525921
rect 331054 525865 331122 525921
rect 331178 525865 361718 525921
rect 361774 525865 361842 525921
rect 361898 525865 392438 525921
rect 392494 525865 392562 525921
rect 392618 525865 423158 525921
rect 423214 525865 423282 525921
rect 423338 525865 453878 525921
rect 453934 525865 454002 525921
rect 454058 525865 484598 525921
rect 484654 525865 484722 525921
rect 484778 525865 515318 525921
rect 515374 525865 515442 525921
rect 515498 525865 546038 525921
rect 546094 525865 546162 525921
rect 546218 525865 597980 525921
rect -1916 525826 597980 525865
rect -1916 514350 597980 514446
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 6970 514350
rect 7026 514294 7094 514350
rect 7150 514294 7218 514350
rect 7274 514294 7342 514350
rect 7398 514294 24970 514350
rect 25026 514294 25094 514350
rect 25150 514294 25218 514350
rect 25274 514294 25342 514350
rect 25398 514294 42970 514350
rect 43026 514294 43094 514350
rect 43150 514294 43218 514350
rect 43274 514294 43342 514350
rect 43398 514294 60970 514350
rect 61026 514294 61094 514350
rect 61150 514294 61218 514350
rect 61274 514294 61342 514350
rect 61398 514294 69878 514350
rect 69934 514294 70002 514350
rect 70058 514294 78970 514350
rect 79026 514294 79094 514350
rect 79150 514294 79218 514350
rect 79274 514294 79342 514350
rect 79398 514294 96970 514350
rect 97026 514294 97094 514350
rect 97150 514294 97218 514350
rect 97274 514294 97342 514350
rect 97398 514294 100598 514350
rect 100654 514294 100722 514350
rect 100778 514294 131318 514350
rect 131374 514294 131442 514350
rect 131498 514294 162038 514350
rect 162094 514294 162162 514350
rect 162218 514294 192758 514350
rect 192814 514294 192882 514350
rect 192938 514294 223478 514350
rect 223534 514294 223602 514350
rect 223658 514294 254198 514350
rect 254254 514294 254322 514350
rect 254378 514294 284918 514350
rect 284974 514294 285042 514350
rect 285098 514294 315638 514350
rect 315694 514294 315762 514350
rect 315818 514294 346358 514350
rect 346414 514294 346482 514350
rect 346538 514294 377078 514350
rect 377134 514294 377202 514350
rect 377258 514294 407798 514350
rect 407854 514294 407922 514350
rect 407978 514294 438518 514350
rect 438574 514294 438642 514350
rect 438698 514294 469238 514350
rect 469294 514294 469362 514350
rect 469418 514294 499958 514350
rect 500014 514294 500082 514350
rect 500138 514294 530678 514350
rect 530734 514294 530802 514350
rect 530858 514294 564970 514350
rect 565026 514294 565094 514350
rect 565150 514294 565218 514350
rect 565274 514294 565342 514350
rect 565398 514294 582970 514350
rect 583026 514294 583094 514350
rect 583150 514294 583218 514350
rect 583274 514294 583342 514350
rect 583398 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect -1916 514226 597980 514294
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 6970 514226
rect 7026 514170 7094 514226
rect 7150 514170 7218 514226
rect 7274 514170 7342 514226
rect 7398 514170 24970 514226
rect 25026 514170 25094 514226
rect 25150 514170 25218 514226
rect 25274 514170 25342 514226
rect 25398 514170 42970 514226
rect 43026 514170 43094 514226
rect 43150 514170 43218 514226
rect 43274 514170 43342 514226
rect 43398 514170 60970 514226
rect 61026 514170 61094 514226
rect 61150 514170 61218 514226
rect 61274 514170 61342 514226
rect 61398 514170 69878 514226
rect 69934 514170 70002 514226
rect 70058 514170 78970 514226
rect 79026 514170 79094 514226
rect 79150 514170 79218 514226
rect 79274 514170 79342 514226
rect 79398 514170 96970 514226
rect 97026 514170 97094 514226
rect 97150 514170 97218 514226
rect 97274 514170 97342 514226
rect 97398 514170 100598 514226
rect 100654 514170 100722 514226
rect 100778 514170 131318 514226
rect 131374 514170 131442 514226
rect 131498 514170 162038 514226
rect 162094 514170 162162 514226
rect 162218 514170 192758 514226
rect 192814 514170 192882 514226
rect 192938 514170 223478 514226
rect 223534 514170 223602 514226
rect 223658 514170 254198 514226
rect 254254 514170 254322 514226
rect 254378 514170 284918 514226
rect 284974 514170 285042 514226
rect 285098 514170 315638 514226
rect 315694 514170 315762 514226
rect 315818 514170 346358 514226
rect 346414 514170 346482 514226
rect 346538 514170 377078 514226
rect 377134 514170 377202 514226
rect 377258 514170 407798 514226
rect 407854 514170 407922 514226
rect 407978 514170 438518 514226
rect 438574 514170 438642 514226
rect 438698 514170 469238 514226
rect 469294 514170 469362 514226
rect 469418 514170 499958 514226
rect 500014 514170 500082 514226
rect 500138 514170 530678 514226
rect 530734 514170 530802 514226
rect 530858 514170 564970 514226
rect 565026 514170 565094 514226
rect 565150 514170 565218 514226
rect 565274 514170 565342 514226
rect 565398 514170 582970 514226
rect 583026 514170 583094 514226
rect 583150 514170 583218 514226
rect 583274 514170 583342 514226
rect 583398 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect -1916 514102 597980 514170
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 6970 514102
rect 7026 514046 7094 514102
rect 7150 514046 7218 514102
rect 7274 514046 7342 514102
rect 7398 514046 24970 514102
rect 25026 514046 25094 514102
rect 25150 514046 25218 514102
rect 25274 514046 25342 514102
rect 25398 514046 42970 514102
rect 43026 514046 43094 514102
rect 43150 514046 43218 514102
rect 43274 514046 43342 514102
rect 43398 514046 60970 514102
rect 61026 514046 61094 514102
rect 61150 514046 61218 514102
rect 61274 514046 61342 514102
rect 61398 514046 69878 514102
rect 69934 514046 70002 514102
rect 70058 514046 78970 514102
rect 79026 514046 79094 514102
rect 79150 514046 79218 514102
rect 79274 514046 79342 514102
rect 79398 514046 96970 514102
rect 97026 514046 97094 514102
rect 97150 514046 97218 514102
rect 97274 514046 97342 514102
rect 97398 514046 100598 514102
rect 100654 514046 100722 514102
rect 100778 514046 131318 514102
rect 131374 514046 131442 514102
rect 131498 514046 162038 514102
rect 162094 514046 162162 514102
rect 162218 514046 192758 514102
rect 192814 514046 192882 514102
rect 192938 514046 223478 514102
rect 223534 514046 223602 514102
rect 223658 514046 254198 514102
rect 254254 514046 254322 514102
rect 254378 514046 284918 514102
rect 284974 514046 285042 514102
rect 285098 514046 315638 514102
rect 315694 514046 315762 514102
rect 315818 514046 346358 514102
rect 346414 514046 346482 514102
rect 346538 514046 377078 514102
rect 377134 514046 377202 514102
rect 377258 514046 407798 514102
rect 407854 514046 407922 514102
rect 407978 514046 438518 514102
rect 438574 514046 438642 514102
rect 438698 514046 469238 514102
rect 469294 514046 469362 514102
rect 469418 514046 499958 514102
rect 500014 514046 500082 514102
rect 500138 514046 530678 514102
rect 530734 514046 530802 514102
rect 530858 514046 564970 514102
rect 565026 514046 565094 514102
rect 565150 514046 565218 514102
rect 565274 514046 565342 514102
rect 565398 514046 582970 514102
rect 583026 514046 583094 514102
rect 583150 514046 583218 514102
rect 583274 514046 583342 514102
rect 583398 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect -1916 513978 597980 514046
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 6970 513978
rect 7026 513922 7094 513978
rect 7150 513922 7218 513978
rect 7274 513922 7342 513978
rect 7398 513922 24970 513978
rect 25026 513922 25094 513978
rect 25150 513922 25218 513978
rect 25274 513922 25342 513978
rect 25398 513922 42970 513978
rect 43026 513922 43094 513978
rect 43150 513922 43218 513978
rect 43274 513922 43342 513978
rect 43398 513922 60970 513978
rect 61026 513922 61094 513978
rect 61150 513922 61218 513978
rect 61274 513922 61342 513978
rect 61398 513922 69878 513978
rect 69934 513922 70002 513978
rect 70058 513922 78970 513978
rect 79026 513922 79094 513978
rect 79150 513922 79218 513978
rect 79274 513922 79342 513978
rect 79398 513922 96970 513978
rect 97026 513922 97094 513978
rect 97150 513922 97218 513978
rect 97274 513922 97342 513978
rect 97398 513922 100598 513978
rect 100654 513922 100722 513978
rect 100778 513922 131318 513978
rect 131374 513922 131442 513978
rect 131498 513922 162038 513978
rect 162094 513922 162162 513978
rect 162218 513922 192758 513978
rect 192814 513922 192882 513978
rect 192938 513922 223478 513978
rect 223534 513922 223602 513978
rect 223658 513922 254198 513978
rect 254254 513922 254322 513978
rect 254378 513922 284918 513978
rect 284974 513922 285042 513978
rect 285098 513922 315638 513978
rect 315694 513922 315762 513978
rect 315818 513922 346358 513978
rect 346414 513922 346482 513978
rect 346538 513922 377078 513978
rect 377134 513922 377202 513978
rect 377258 513922 407798 513978
rect 407854 513922 407922 513978
rect 407978 513922 438518 513978
rect 438574 513922 438642 513978
rect 438698 513922 469238 513978
rect 469294 513922 469362 513978
rect 469418 513922 499958 513978
rect 500014 513922 500082 513978
rect 500138 513922 530678 513978
rect 530734 513922 530802 513978
rect 530858 513922 564970 513978
rect 565026 513922 565094 513978
rect 565150 513922 565218 513978
rect 565274 513922 565342 513978
rect 565398 513922 582970 513978
rect 583026 513922 583094 513978
rect 583150 513922 583218 513978
rect 583274 513922 583342 513978
rect 583398 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect -1916 513826 597980 513922
rect -1916 508350 597980 508446
rect -1916 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 3250 508350
rect 3306 508294 3374 508350
rect 3430 508294 3498 508350
rect 3554 508294 3622 508350
rect 3678 508294 21250 508350
rect 21306 508294 21374 508350
rect 21430 508294 21498 508350
rect 21554 508294 21622 508350
rect 21678 508294 39250 508350
rect 39306 508294 39374 508350
rect 39430 508294 39498 508350
rect 39554 508294 39622 508350
rect 39678 508294 54518 508350
rect 54574 508294 54642 508350
rect 54698 508294 57250 508350
rect 57306 508294 57374 508350
rect 57430 508294 57498 508350
rect 57554 508294 57622 508350
rect 57678 508294 75250 508350
rect 75306 508294 75374 508350
rect 75430 508294 75498 508350
rect 75554 508294 75622 508350
rect 75678 508294 85238 508350
rect 85294 508294 85362 508350
rect 85418 508294 93250 508350
rect 93306 508294 93374 508350
rect 93430 508294 93498 508350
rect 93554 508294 93622 508350
rect 93678 508294 111250 508350
rect 111306 508294 111374 508350
rect 111430 508294 111498 508350
rect 111554 508294 111622 508350
rect 111678 508294 115958 508350
rect 116014 508294 116082 508350
rect 116138 508294 146678 508350
rect 146734 508294 146802 508350
rect 146858 508294 177398 508350
rect 177454 508294 177522 508350
rect 177578 508294 208118 508350
rect 208174 508294 208242 508350
rect 208298 508294 238838 508350
rect 238894 508294 238962 508350
rect 239018 508294 269558 508350
rect 269614 508294 269682 508350
rect 269738 508294 300278 508350
rect 300334 508294 300402 508350
rect 300458 508294 330998 508350
rect 331054 508294 331122 508350
rect 331178 508294 361718 508350
rect 361774 508294 361842 508350
rect 361898 508294 392438 508350
rect 392494 508294 392562 508350
rect 392618 508294 423158 508350
rect 423214 508294 423282 508350
rect 423338 508294 453878 508350
rect 453934 508294 454002 508350
rect 454058 508294 484598 508350
rect 484654 508294 484722 508350
rect 484778 508294 515318 508350
rect 515374 508294 515442 508350
rect 515498 508294 546038 508350
rect 546094 508294 546162 508350
rect 546218 508294 561250 508350
rect 561306 508294 561374 508350
rect 561430 508294 561498 508350
rect 561554 508294 561622 508350
rect 561678 508294 579250 508350
rect 579306 508294 579374 508350
rect 579430 508294 579498 508350
rect 579554 508294 579622 508350
rect 579678 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597980 508350
rect -1916 508226 597980 508294
rect -1916 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 3250 508226
rect 3306 508170 3374 508226
rect 3430 508170 3498 508226
rect 3554 508170 3622 508226
rect 3678 508170 21250 508226
rect 21306 508170 21374 508226
rect 21430 508170 21498 508226
rect 21554 508170 21622 508226
rect 21678 508170 39250 508226
rect 39306 508170 39374 508226
rect 39430 508170 39498 508226
rect 39554 508170 39622 508226
rect 39678 508170 54518 508226
rect 54574 508170 54642 508226
rect 54698 508170 57250 508226
rect 57306 508170 57374 508226
rect 57430 508170 57498 508226
rect 57554 508170 57622 508226
rect 57678 508170 75250 508226
rect 75306 508170 75374 508226
rect 75430 508170 75498 508226
rect 75554 508170 75622 508226
rect 75678 508170 85238 508226
rect 85294 508170 85362 508226
rect 85418 508170 93250 508226
rect 93306 508170 93374 508226
rect 93430 508170 93498 508226
rect 93554 508170 93622 508226
rect 93678 508170 111250 508226
rect 111306 508170 111374 508226
rect 111430 508170 111498 508226
rect 111554 508170 111622 508226
rect 111678 508170 115958 508226
rect 116014 508170 116082 508226
rect 116138 508170 146678 508226
rect 146734 508170 146802 508226
rect 146858 508170 177398 508226
rect 177454 508170 177522 508226
rect 177578 508170 208118 508226
rect 208174 508170 208242 508226
rect 208298 508170 238838 508226
rect 238894 508170 238962 508226
rect 239018 508170 269558 508226
rect 269614 508170 269682 508226
rect 269738 508170 300278 508226
rect 300334 508170 300402 508226
rect 300458 508170 330998 508226
rect 331054 508170 331122 508226
rect 331178 508170 361718 508226
rect 361774 508170 361842 508226
rect 361898 508170 392438 508226
rect 392494 508170 392562 508226
rect 392618 508170 423158 508226
rect 423214 508170 423282 508226
rect 423338 508170 453878 508226
rect 453934 508170 454002 508226
rect 454058 508170 484598 508226
rect 484654 508170 484722 508226
rect 484778 508170 515318 508226
rect 515374 508170 515442 508226
rect 515498 508170 546038 508226
rect 546094 508170 546162 508226
rect 546218 508170 561250 508226
rect 561306 508170 561374 508226
rect 561430 508170 561498 508226
rect 561554 508170 561622 508226
rect 561678 508170 579250 508226
rect 579306 508170 579374 508226
rect 579430 508170 579498 508226
rect 579554 508170 579622 508226
rect 579678 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597980 508226
rect -1916 508102 597980 508170
rect -1916 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 3250 508102
rect 3306 508046 3374 508102
rect 3430 508046 3498 508102
rect 3554 508046 3622 508102
rect 3678 508046 21250 508102
rect 21306 508046 21374 508102
rect 21430 508046 21498 508102
rect 21554 508046 21622 508102
rect 21678 508046 39250 508102
rect 39306 508046 39374 508102
rect 39430 508046 39498 508102
rect 39554 508046 39622 508102
rect 39678 508046 54518 508102
rect 54574 508046 54642 508102
rect 54698 508046 57250 508102
rect 57306 508046 57374 508102
rect 57430 508046 57498 508102
rect 57554 508046 57622 508102
rect 57678 508046 75250 508102
rect 75306 508046 75374 508102
rect 75430 508046 75498 508102
rect 75554 508046 75622 508102
rect 75678 508046 85238 508102
rect 85294 508046 85362 508102
rect 85418 508046 93250 508102
rect 93306 508046 93374 508102
rect 93430 508046 93498 508102
rect 93554 508046 93622 508102
rect 93678 508046 111250 508102
rect 111306 508046 111374 508102
rect 111430 508046 111498 508102
rect 111554 508046 111622 508102
rect 111678 508046 115958 508102
rect 116014 508046 116082 508102
rect 116138 508046 146678 508102
rect 146734 508046 146802 508102
rect 146858 508046 177398 508102
rect 177454 508046 177522 508102
rect 177578 508046 208118 508102
rect 208174 508046 208242 508102
rect 208298 508046 238838 508102
rect 238894 508046 238962 508102
rect 239018 508046 269558 508102
rect 269614 508046 269682 508102
rect 269738 508046 300278 508102
rect 300334 508046 300402 508102
rect 300458 508046 330998 508102
rect 331054 508046 331122 508102
rect 331178 508046 361718 508102
rect 361774 508046 361842 508102
rect 361898 508046 392438 508102
rect 392494 508046 392562 508102
rect 392618 508046 423158 508102
rect 423214 508046 423282 508102
rect 423338 508046 453878 508102
rect 453934 508046 454002 508102
rect 454058 508046 484598 508102
rect 484654 508046 484722 508102
rect 484778 508046 515318 508102
rect 515374 508046 515442 508102
rect 515498 508046 546038 508102
rect 546094 508046 546162 508102
rect 546218 508046 561250 508102
rect 561306 508046 561374 508102
rect 561430 508046 561498 508102
rect 561554 508046 561622 508102
rect 561678 508046 579250 508102
rect 579306 508046 579374 508102
rect 579430 508046 579498 508102
rect 579554 508046 579622 508102
rect 579678 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597980 508102
rect -1916 507978 597980 508046
rect -1916 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 3250 507978
rect 3306 507922 3374 507978
rect 3430 507922 3498 507978
rect 3554 507922 3622 507978
rect 3678 507922 21250 507978
rect 21306 507922 21374 507978
rect 21430 507922 21498 507978
rect 21554 507922 21622 507978
rect 21678 507922 39250 507978
rect 39306 507922 39374 507978
rect 39430 507922 39498 507978
rect 39554 507922 39622 507978
rect 39678 507922 54518 507978
rect 54574 507922 54642 507978
rect 54698 507922 57250 507978
rect 57306 507922 57374 507978
rect 57430 507922 57498 507978
rect 57554 507922 57622 507978
rect 57678 507922 75250 507978
rect 75306 507922 75374 507978
rect 75430 507922 75498 507978
rect 75554 507922 75622 507978
rect 75678 507922 85238 507978
rect 85294 507922 85362 507978
rect 85418 507922 93250 507978
rect 93306 507922 93374 507978
rect 93430 507922 93498 507978
rect 93554 507922 93622 507978
rect 93678 507922 111250 507978
rect 111306 507922 111374 507978
rect 111430 507922 111498 507978
rect 111554 507922 111622 507978
rect 111678 507922 115958 507978
rect 116014 507922 116082 507978
rect 116138 507922 146678 507978
rect 146734 507922 146802 507978
rect 146858 507922 177398 507978
rect 177454 507922 177522 507978
rect 177578 507922 208118 507978
rect 208174 507922 208242 507978
rect 208298 507922 238838 507978
rect 238894 507922 238962 507978
rect 239018 507922 269558 507978
rect 269614 507922 269682 507978
rect 269738 507922 300278 507978
rect 300334 507922 300402 507978
rect 300458 507922 330998 507978
rect 331054 507922 331122 507978
rect 331178 507922 361718 507978
rect 361774 507922 361842 507978
rect 361898 507922 392438 507978
rect 392494 507922 392562 507978
rect 392618 507922 423158 507978
rect 423214 507922 423282 507978
rect 423338 507922 453878 507978
rect 453934 507922 454002 507978
rect 454058 507922 484598 507978
rect 484654 507922 484722 507978
rect 484778 507922 515318 507978
rect 515374 507922 515442 507978
rect 515498 507922 546038 507978
rect 546094 507922 546162 507978
rect 546218 507922 561250 507978
rect 561306 507922 561374 507978
rect 561430 507922 561498 507978
rect 561554 507922 561622 507978
rect 561678 507922 579250 507978
rect 579306 507922 579374 507978
rect 579430 507922 579498 507978
rect 579554 507922 579622 507978
rect 579678 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597980 507978
rect -1916 507826 597980 507922
rect -1916 496350 597980 496446
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 6970 496350
rect 7026 496294 7094 496350
rect 7150 496294 7218 496350
rect 7274 496294 7342 496350
rect 7398 496294 24970 496350
rect 25026 496294 25094 496350
rect 25150 496294 25218 496350
rect 25274 496294 25342 496350
rect 25398 496294 42970 496350
rect 43026 496294 43094 496350
rect 43150 496294 43218 496350
rect 43274 496294 43342 496350
rect 43398 496294 60970 496350
rect 61026 496294 61094 496350
rect 61150 496294 61218 496350
rect 61274 496294 61342 496350
rect 61398 496294 69878 496350
rect 69934 496294 70002 496350
rect 70058 496294 78970 496350
rect 79026 496294 79094 496350
rect 79150 496294 79218 496350
rect 79274 496294 79342 496350
rect 79398 496294 96970 496350
rect 97026 496294 97094 496350
rect 97150 496294 97218 496350
rect 97274 496294 97342 496350
rect 97398 496294 100598 496350
rect 100654 496294 100722 496350
rect 100778 496294 131318 496350
rect 131374 496294 131442 496350
rect 131498 496294 162038 496350
rect 162094 496294 162162 496350
rect 162218 496294 192758 496350
rect 192814 496294 192882 496350
rect 192938 496294 223478 496350
rect 223534 496294 223602 496350
rect 223658 496294 254198 496350
rect 254254 496294 254322 496350
rect 254378 496294 284918 496350
rect 284974 496294 285042 496350
rect 285098 496294 315638 496350
rect 315694 496294 315762 496350
rect 315818 496294 346358 496350
rect 346414 496294 346482 496350
rect 346538 496294 377078 496350
rect 377134 496294 377202 496350
rect 377258 496294 407798 496350
rect 407854 496294 407922 496350
rect 407978 496294 438518 496350
rect 438574 496294 438642 496350
rect 438698 496294 469238 496350
rect 469294 496294 469362 496350
rect 469418 496294 499958 496350
rect 500014 496294 500082 496350
rect 500138 496294 530678 496350
rect 530734 496294 530802 496350
rect 530858 496294 564970 496350
rect 565026 496294 565094 496350
rect 565150 496294 565218 496350
rect 565274 496294 565342 496350
rect 565398 496294 582970 496350
rect 583026 496294 583094 496350
rect 583150 496294 583218 496350
rect 583274 496294 583342 496350
rect 583398 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect -1916 496226 597980 496294
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 6970 496226
rect 7026 496170 7094 496226
rect 7150 496170 7218 496226
rect 7274 496170 7342 496226
rect 7398 496170 24970 496226
rect 25026 496170 25094 496226
rect 25150 496170 25218 496226
rect 25274 496170 25342 496226
rect 25398 496170 42970 496226
rect 43026 496170 43094 496226
rect 43150 496170 43218 496226
rect 43274 496170 43342 496226
rect 43398 496170 60970 496226
rect 61026 496170 61094 496226
rect 61150 496170 61218 496226
rect 61274 496170 61342 496226
rect 61398 496170 69878 496226
rect 69934 496170 70002 496226
rect 70058 496170 78970 496226
rect 79026 496170 79094 496226
rect 79150 496170 79218 496226
rect 79274 496170 79342 496226
rect 79398 496170 96970 496226
rect 97026 496170 97094 496226
rect 97150 496170 97218 496226
rect 97274 496170 97342 496226
rect 97398 496170 100598 496226
rect 100654 496170 100722 496226
rect 100778 496170 131318 496226
rect 131374 496170 131442 496226
rect 131498 496170 162038 496226
rect 162094 496170 162162 496226
rect 162218 496170 192758 496226
rect 192814 496170 192882 496226
rect 192938 496170 223478 496226
rect 223534 496170 223602 496226
rect 223658 496170 254198 496226
rect 254254 496170 254322 496226
rect 254378 496170 284918 496226
rect 284974 496170 285042 496226
rect 285098 496170 315638 496226
rect 315694 496170 315762 496226
rect 315818 496170 346358 496226
rect 346414 496170 346482 496226
rect 346538 496170 377078 496226
rect 377134 496170 377202 496226
rect 377258 496170 407798 496226
rect 407854 496170 407922 496226
rect 407978 496170 438518 496226
rect 438574 496170 438642 496226
rect 438698 496170 469238 496226
rect 469294 496170 469362 496226
rect 469418 496170 499958 496226
rect 500014 496170 500082 496226
rect 500138 496170 530678 496226
rect 530734 496170 530802 496226
rect 530858 496170 564970 496226
rect 565026 496170 565094 496226
rect 565150 496170 565218 496226
rect 565274 496170 565342 496226
rect 565398 496170 582970 496226
rect 583026 496170 583094 496226
rect 583150 496170 583218 496226
rect 583274 496170 583342 496226
rect 583398 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect -1916 496102 597980 496170
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 6970 496102
rect 7026 496046 7094 496102
rect 7150 496046 7218 496102
rect 7274 496046 7342 496102
rect 7398 496046 24970 496102
rect 25026 496046 25094 496102
rect 25150 496046 25218 496102
rect 25274 496046 25342 496102
rect 25398 496046 42970 496102
rect 43026 496046 43094 496102
rect 43150 496046 43218 496102
rect 43274 496046 43342 496102
rect 43398 496046 60970 496102
rect 61026 496046 61094 496102
rect 61150 496046 61218 496102
rect 61274 496046 61342 496102
rect 61398 496046 69878 496102
rect 69934 496046 70002 496102
rect 70058 496046 78970 496102
rect 79026 496046 79094 496102
rect 79150 496046 79218 496102
rect 79274 496046 79342 496102
rect 79398 496046 96970 496102
rect 97026 496046 97094 496102
rect 97150 496046 97218 496102
rect 97274 496046 97342 496102
rect 97398 496046 100598 496102
rect 100654 496046 100722 496102
rect 100778 496046 131318 496102
rect 131374 496046 131442 496102
rect 131498 496046 162038 496102
rect 162094 496046 162162 496102
rect 162218 496046 192758 496102
rect 192814 496046 192882 496102
rect 192938 496046 223478 496102
rect 223534 496046 223602 496102
rect 223658 496046 254198 496102
rect 254254 496046 254322 496102
rect 254378 496046 284918 496102
rect 284974 496046 285042 496102
rect 285098 496046 315638 496102
rect 315694 496046 315762 496102
rect 315818 496046 346358 496102
rect 346414 496046 346482 496102
rect 346538 496046 377078 496102
rect 377134 496046 377202 496102
rect 377258 496046 407798 496102
rect 407854 496046 407922 496102
rect 407978 496046 438518 496102
rect 438574 496046 438642 496102
rect 438698 496046 469238 496102
rect 469294 496046 469362 496102
rect 469418 496046 499958 496102
rect 500014 496046 500082 496102
rect 500138 496046 530678 496102
rect 530734 496046 530802 496102
rect 530858 496046 564970 496102
rect 565026 496046 565094 496102
rect 565150 496046 565218 496102
rect 565274 496046 565342 496102
rect 565398 496046 582970 496102
rect 583026 496046 583094 496102
rect 583150 496046 583218 496102
rect 583274 496046 583342 496102
rect 583398 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect -1916 495978 597980 496046
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 6970 495978
rect 7026 495922 7094 495978
rect 7150 495922 7218 495978
rect 7274 495922 7342 495978
rect 7398 495922 24970 495978
rect 25026 495922 25094 495978
rect 25150 495922 25218 495978
rect 25274 495922 25342 495978
rect 25398 495922 42970 495978
rect 43026 495922 43094 495978
rect 43150 495922 43218 495978
rect 43274 495922 43342 495978
rect 43398 495922 60970 495978
rect 61026 495922 61094 495978
rect 61150 495922 61218 495978
rect 61274 495922 61342 495978
rect 61398 495922 69878 495978
rect 69934 495922 70002 495978
rect 70058 495922 78970 495978
rect 79026 495922 79094 495978
rect 79150 495922 79218 495978
rect 79274 495922 79342 495978
rect 79398 495922 96970 495978
rect 97026 495922 97094 495978
rect 97150 495922 97218 495978
rect 97274 495922 97342 495978
rect 97398 495922 100598 495978
rect 100654 495922 100722 495978
rect 100778 495922 131318 495978
rect 131374 495922 131442 495978
rect 131498 495922 162038 495978
rect 162094 495922 162162 495978
rect 162218 495922 192758 495978
rect 192814 495922 192882 495978
rect 192938 495922 223478 495978
rect 223534 495922 223602 495978
rect 223658 495922 254198 495978
rect 254254 495922 254322 495978
rect 254378 495922 284918 495978
rect 284974 495922 285042 495978
rect 285098 495922 315638 495978
rect 315694 495922 315762 495978
rect 315818 495922 346358 495978
rect 346414 495922 346482 495978
rect 346538 495922 377078 495978
rect 377134 495922 377202 495978
rect 377258 495922 407798 495978
rect 407854 495922 407922 495978
rect 407978 495922 438518 495978
rect 438574 495922 438642 495978
rect 438698 495922 469238 495978
rect 469294 495922 469362 495978
rect 469418 495922 499958 495978
rect 500014 495922 500082 495978
rect 500138 495922 530678 495978
rect 530734 495922 530802 495978
rect 530858 495922 564970 495978
rect 565026 495922 565094 495978
rect 565150 495922 565218 495978
rect 565274 495922 565342 495978
rect 565398 495922 582970 495978
rect 583026 495922 583094 495978
rect 583150 495922 583218 495978
rect 583274 495922 583342 495978
rect 583398 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect -1916 495826 597980 495922
rect -1916 490350 597980 490446
rect -1916 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 3250 490350
rect 3306 490294 3374 490350
rect 3430 490294 3498 490350
rect 3554 490294 3622 490350
rect 3678 490294 21250 490350
rect 21306 490294 21374 490350
rect 21430 490294 21498 490350
rect 21554 490294 21622 490350
rect 21678 490294 39250 490350
rect 39306 490294 39374 490350
rect 39430 490294 39498 490350
rect 39554 490294 39622 490350
rect 39678 490294 54518 490350
rect 54574 490294 54642 490350
rect 54698 490294 57250 490350
rect 57306 490294 57374 490350
rect 57430 490294 57498 490350
rect 57554 490294 57622 490350
rect 57678 490294 75250 490350
rect 75306 490294 75374 490350
rect 75430 490294 75498 490350
rect 75554 490294 75622 490350
rect 75678 490294 85238 490350
rect 85294 490294 85362 490350
rect 85418 490294 93250 490350
rect 93306 490294 93374 490350
rect 93430 490294 93498 490350
rect 93554 490294 93622 490350
rect 93678 490294 111250 490350
rect 111306 490294 111374 490350
rect 111430 490294 111498 490350
rect 111554 490294 111622 490350
rect 111678 490294 115958 490350
rect 116014 490294 116082 490350
rect 116138 490294 146678 490350
rect 146734 490294 146802 490350
rect 146858 490294 177398 490350
rect 177454 490294 177522 490350
rect 177578 490294 208118 490350
rect 208174 490294 208242 490350
rect 208298 490294 238838 490350
rect 238894 490294 238962 490350
rect 239018 490294 269558 490350
rect 269614 490294 269682 490350
rect 269738 490294 300278 490350
rect 300334 490294 300402 490350
rect 300458 490294 330998 490350
rect 331054 490294 331122 490350
rect 331178 490294 361718 490350
rect 361774 490294 361842 490350
rect 361898 490294 392438 490350
rect 392494 490294 392562 490350
rect 392618 490294 423158 490350
rect 423214 490294 423282 490350
rect 423338 490294 453878 490350
rect 453934 490294 454002 490350
rect 454058 490294 484598 490350
rect 484654 490294 484722 490350
rect 484778 490294 515318 490350
rect 515374 490294 515442 490350
rect 515498 490294 546038 490350
rect 546094 490294 546162 490350
rect 546218 490294 561250 490350
rect 561306 490294 561374 490350
rect 561430 490294 561498 490350
rect 561554 490294 561622 490350
rect 561678 490294 579250 490350
rect 579306 490294 579374 490350
rect 579430 490294 579498 490350
rect 579554 490294 579622 490350
rect 579678 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597980 490350
rect -1916 490226 597980 490294
rect -1916 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 3250 490226
rect 3306 490170 3374 490226
rect 3430 490170 3498 490226
rect 3554 490170 3622 490226
rect 3678 490170 21250 490226
rect 21306 490170 21374 490226
rect 21430 490170 21498 490226
rect 21554 490170 21622 490226
rect 21678 490170 39250 490226
rect 39306 490170 39374 490226
rect 39430 490170 39498 490226
rect 39554 490170 39622 490226
rect 39678 490170 54518 490226
rect 54574 490170 54642 490226
rect 54698 490170 57250 490226
rect 57306 490170 57374 490226
rect 57430 490170 57498 490226
rect 57554 490170 57622 490226
rect 57678 490170 75250 490226
rect 75306 490170 75374 490226
rect 75430 490170 75498 490226
rect 75554 490170 75622 490226
rect 75678 490170 85238 490226
rect 85294 490170 85362 490226
rect 85418 490170 93250 490226
rect 93306 490170 93374 490226
rect 93430 490170 93498 490226
rect 93554 490170 93622 490226
rect 93678 490170 111250 490226
rect 111306 490170 111374 490226
rect 111430 490170 111498 490226
rect 111554 490170 111622 490226
rect 111678 490170 115958 490226
rect 116014 490170 116082 490226
rect 116138 490170 146678 490226
rect 146734 490170 146802 490226
rect 146858 490170 177398 490226
rect 177454 490170 177522 490226
rect 177578 490170 208118 490226
rect 208174 490170 208242 490226
rect 208298 490170 238838 490226
rect 238894 490170 238962 490226
rect 239018 490170 269558 490226
rect 269614 490170 269682 490226
rect 269738 490170 300278 490226
rect 300334 490170 300402 490226
rect 300458 490170 330998 490226
rect 331054 490170 331122 490226
rect 331178 490170 361718 490226
rect 361774 490170 361842 490226
rect 361898 490170 392438 490226
rect 392494 490170 392562 490226
rect 392618 490170 423158 490226
rect 423214 490170 423282 490226
rect 423338 490170 453878 490226
rect 453934 490170 454002 490226
rect 454058 490170 484598 490226
rect 484654 490170 484722 490226
rect 484778 490170 515318 490226
rect 515374 490170 515442 490226
rect 515498 490170 546038 490226
rect 546094 490170 546162 490226
rect 546218 490170 561250 490226
rect 561306 490170 561374 490226
rect 561430 490170 561498 490226
rect 561554 490170 561622 490226
rect 561678 490170 579250 490226
rect 579306 490170 579374 490226
rect 579430 490170 579498 490226
rect 579554 490170 579622 490226
rect 579678 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597980 490226
rect -1916 490102 597980 490170
rect -1916 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 3250 490102
rect 3306 490046 3374 490102
rect 3430 490046 3498 490102
rect 3554 490046 3622 490102
rect 3678 490046 21250 490102
rect 21306 490046 21374 490102
rect 21430 490046 21498 490102
rect 21554 490046 21622 490102
rect 21678 490046 39250 490102
rect 39306 490046 39374 490102
rect 39430 490046 39498 490102
rect 39554 490046 39622 490102
rect 39678 490046 54518 490102
rect 54574 490046 54642 490102
rect 54698 490046 57250 490102
rect 57306 490046 57374 490102
rect 57430 490046 57498 490102
rect 57554 490046 57622 490102
rect 57678 490046 75250 490102
rect 75306 490046 75374 490102
rect 75430 490046 75498 490102
rect 75554 490046 75622 490102
rect 75678 490046 85238 490102
rect 85294 490046 85362 490102
rect 85418 490046 93250 490102
rect 93306 490046 93374 490102
rect 93430 490046 93498 490102
rect 93554 490046 93622 490102
rect 93678 490046 111250 490102
rect 111306 490046 111374 490102
rect 111430 490046 111498 490102
rect 111554 490046 111622 490102
rect 111678 490046 115958 490102
rect 116014 490046 116082 490102
rect 116138 490046 146678 490102
rect 146734 490046 146802 490102
rect 146858 490046 177398 490102
rect 177454 490046 177522 490102
rect 177578 490046 208118 490102
rect 208174 490046 208242 490102
rect 208298 490046 238838 490102
rect 238894 490046 238962 490102
rect 239018 490046 269558 490102
rect 269614 490046 269682 490102
rect 269738 490046 300278 490102
rect 300334 490046 300402 490102
rect 300458 490046 330998 490102
rect 331054 490046 331122 490102
rect 331178 490046 361718 490102
rect 361774 490046 361842 490102
rect 361898 490046 392438 490102
rect 392494 490046 392562 490102
rect 392618 490046 423158 490102
rect 423214 490046 423282 490102
rect 423338 490046 453878 490102
rect 453934 490046 454002 490102
rect 454058 490046 484598 490102
rect 484654 490046 484722 490102
rect 484778 490046 515318 490102
rect 515374 490046 515442 490102
rect 515498 490046 546038 490102
rect 546094 490046 546162 490102
rect 546218 490046 561250 490102
rect 561306 490046 561374 490102
rect 561430 490046 561498 490102
rect 561554 490046 561622 490102
rect 561678 490046 579250 490102
rect 579306 490046 579374 490102
rect 579430 490046 579498 490102
rect 579554 490046 579622 490102
rect 579678 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597980 490102
rect -1916 489978 597980 490046
rect -1916 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 3250 489978
rect 3306 489922 3374 489978
rect 3430 489922 3498 489978
rect 3554 489922 3622 489978
rect 3678 489922 21250 489978
rect 21306 489922 21374 489978
rect 21430 489922 21498 489978
rect 21554 489922 21622 489978
rect 21678 489922 39250 489978
rect 39306 489922 39374 489978
rect 39430 489922 39498 489978
rect 39554 489922 39622 489978
rect 39678 489922 54518 489978
rect 54574 489922 54642 489978
rect 54698 489922 57250 489978
rect 57306 489922 57374 489978
rect 57430 489922 57498 489978
rect 57554 489922 57622 489978
rect 57678 489922 75250 489978
rect 75306 489922 75374 489978
rect 75430 489922 75498 489978
rect 75554 489922 75622 489978
rect 75678 489922 85238 489978
rect 85294 489922 85362 489978
rect 85418 489922 93250 489978
rect 93306 489922 93374 489978
rect 93430 489922 93498 489978
rect 93554 489922 93622 489978
rect 93678 489922 111250 489978
rect 111306 489922 111374 489978
rect 111430 489922 111498 489978
rect 111554 489922 111622 489978
rect 111678 489922 115958 489978
rect 116014 489922 116082 489978
rect 116138 489922 146678 489978
rect 146734 489922 146802 489978
rect 146858 489922 177398 489978
rect 177454 489922 177522 489978
rect 177578 489922 208118 489978
rect 208174 489922 208242 489978
rect 208298 489922 238838 489978
rect 238894 489922 238962 489978
rect 239018 489922 269558 489978
rect 269614 489922 269682 489978
rect 269738 489922 300278 489978
rect 300334 489922 300402 489978
rect 300458 489922 330998 489978
rect 331054 489922 331122 489978
rect 331178 489922 361718 489978
rect 361774 489922 361842 489978
rect 361898 489922 392438 489978
rect 392494 489922 392562 489978
rect 392618 489922 423158 489978
rect 423214 489922 423282 489978
rect 423338 489922 453878 489978
rect 453934 489922 454002 489978
rect 454058 489922 484598 489978
rect 484654 489922 484722 489978
rect 484778 489922 515318 489978
rect 515374 489922 515442 489978
rect 515498 489922 546038 489978
rect 546094 489922 546162 489978
rect 546218 489922 561250 489978
rect 561306 489922 561374 489978
rect 561430 489922 561498 489978
rect 561554 489922 561622 489978
rect 561678 489922 579250 489978
rect 579306 489922 579374 489978
rect 579430 489922 579498 489978
rect 579554 489922 579622 489978
rect 579678 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597980 489978
rect -1916 489826 597980 489922
rect -1916 478350 597980 478446
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 6970 478350
rect 7026 478294 7094 478350
rect 7150 478294 7218 478350
rect 7274 478294 7342 478350
rect 7398 478294 24970 478350
rect 25026 478294 25094 478350
rect 25150 478294 25218 478350
rect 25274 478294 25342 478350
rect 25398 478294 42970 478350
rect 43026 478294 43094 478350
rect 43150 478294 43218 478350
rect 43274 478294 43342 478350
rect 43398 478294 60970 478350
rect 61026 478294 61094 478350
rect 61150 478294 61218 478350
rect 61274 478294 61342 478350
rect 61398 478294 69878 478350
rect 69934 478294 70002 478350
rect 70058 478294 78970 478350
rect 79026 478294 79094 478350
rect 79150 478294 79218 478350
rect 79274 478294 79342 478350
rect 79398 478294 96970 478350
rect 97026 478294 97094 478350
rect 97150 478294 97218 478350
rect 97274 478294 97342 478350
rect 97398 478294 100598 478350
rect 100654 478294 100722 478350
rect 100778 478294 131318 478350
rect 131374 478294 131442 478350
rect 131498 478294 162038 478350
rect 162094 478294 162162 478350
rect 162218 478294 192758 478350
rect 192814 478294 192882 478350
rect 192938 478294 223478 478350
rect 223534 478294 223602 478350
rect 223658 478294 254198 478350
rect 254254 478294 254322 478350
rect 254378 478294 284918 478350
rect 284974 478294 285042 478350
rect 285098 478294 315638 478350
rect 315694 478294 315762 478350
rect 315818 478294 346358 478350
rect 346414 478294 346482 478350
rect 346538 478294 377078 478350
rect 377134 478294 377202 478350
rect 377258 478294 407798 478350
rect 407854 478294 407922 478350
rect 407978 478294 438518 478350
rect 438574 478294 438642 478350
rect 438698 478294 469238 478350
rect 469294 478294 469362 478350
rect 469418 478294 499958 478350
rect 500014 478294 500082 478350
rect 500138 478294 530678 478350
rect 530734 478294 530802 478350
rect 530858 478294 564970 478350
rect 565026 478294 565094 478350
rect 565150 478294 565218 478350
rect 565274 478294 565342 478350
rect 565398 478294 582970 478350
rect 583026 478294 583094 478350
rect 583150 478294 583218 478350
rect 583274 478294 583342 478350
rect 583398 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect -1916 478226 597980 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 6970 478226
rect 7026 478170 7094 478226
rect 7150 478170 7218 478226
rect 7274 478170 7342 478226
rect 7398 478170 24970 478226
rect 25026 478170 25094 478226
rect 25150 478170 25218 478226
rect 25274 478170 25342 478226
rect 25398 478170 42970 478226
rect 43026 478170 43094 478226
rect 43150 478170 43218 478226
rect 43274 478170 43342 478226
rect 43398 478170 60970 478226
rect 61026 478170 61094 478226
rect 61150 478170 61218 478226
rect 61274 478170 61342 478226
rect 61398 478170 69878 478226
rect 69934 478170 70002 478226
rect 70058 478170 78970 478226
rect 79026 478170 79094 478226
rect 79150 478170 79218 478226
rect 79274 478170 79342 478226
rect 79398 478170 96970 478226
rect 97026 478170 97094 478226
rect 97150 478170 97218 478226
rect 97274 478170 97342 478226
rect 97398 478170 100598 478226
rect 100654 478170 100722 478226
rect 100778 478170 131318 478226
rect 131374 478170 131442 478226
rect 131498 478170 162038 478226
rect 162094 478170 162162 478226
rect 162218 478170 192758 478226
rect 192814 478170 192882 478226
rect 192938 478170 223478 478226
rect 223534 478170 223602 478226
rect 223658 478170 254198 478226
rect 254254 478170 254322 478226
rect 254378 478170 284918 478226
rect 284974 478170 285042 478226
rect 285098 478170 315638 478226
rect 315694 478170 315762 478226
rect 315818 478170 346358 478226
rect 346414 478170 346482 478226
rect 346538 478170 377078 478226
rect 377134 478170 377202 478226
rect 377258 478170 407798 478226
rect 407854 478170 407922 478226
rect 407978 478170 438518 478226
rect 438574 478170 438642 478226
rect 438698 478170 469238 478226
rect 469294 478170 469362 478226
rect 469418 478170 499958 478226
rect 500014 478170 500082 478226
rect 500138 478170 530678 478226
rect 530734 478170 530802 478226
rect 530858 478170 564970 478226
rect 565026 478170 565094 478226
rect 565150 478170 565218 478226
rect 565274 478170 565342 478226
rect 565398 478170 582970 478226
rect 583026 478170 583094 478226
rect 583150 478170 583218 478226
rect 583274 478170 583342 478226
rect 583398 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect -1916 478102 597980 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 6970 478102
rect 7026 478046 7094 478102
rect 7150 478046 7218 478102
rect 7274 478046 7342 478102
rect 7398 478046 24970 478102
rect 25026 478046 25094 478102
rect 25150 478046 25218 478102
rect 25274 478046 25342 478102
rect 25398 478046 42970 478102
rect 43026 478046 43094 478102
rect 43150 478046 43218 478102
rect 43274 478046 43342 478102
rect 43398 478046 60970 478102
rect 61026 478046 61094 478102
rect 61150 478046 61218 478102
rect 61274 478046 61342 478102
rect 61398 478046 69878 478102
rect 69934 478046 70002 478102
rect 70058 478046 78970 478102
rect 79026 478046 79094 478102
rect 79150 478046 79218 478102
rect 79274 478046 79342 478102
rect 79398 478046 96970 478102
rect 97026 478046 97094 478102
rect 97150 478046 97218 478102
rect 97274 478046 97342 478102
rect 97398 478046 100598 478102
rect 100654 478046 100722 478102
rect 100778 478046 131318 478102
rect 131374 478046 131442 478102
rect 131498 478046 162038 478102
rect 162094 478046 162162 478102
rect 162218 478046 192758 478102
rect 192814 478046 192882 478102
rect 192938 478046 223478 478102
rect 223534 478046 223602 478102
rect 223658 478046 254198 478102
rect 254254 478046 254322 478102
rect 254378 478046 284918 478102
rect 284974 478046 285042 478102
rect 285098 478046 315638 478102
rect 315694 478046 315762 478102
rect 315818 478046 346358 478102
rect 346414 478046 346482 478102
rect 346538 478046 377078 478102
rect 377134 478046 377202 478102
rect 377258 478046 407798 478102
rect 407854 478046 407922 478102
rect 407978 478046 438518 478102
rect 438574 478046 438642 478102
rect 438698 478046 469238 478102
rect 469294 478046 469362 478102
rect 469418 478046 499958 478102
rect 500014 478046 500082 478102
rect 500138 478046 530678 478102
rect 530734 478046 530802 478102
rect 530858 478046 564970 478102
rect 565026 478046 565094 478102
rect 565150 478046 565218 478102
rect 565274 478046 565342 478102
rect 565398 478046 582970 478102
rect 583026 478046 583094 478102
rect 583150 478046 583218 478102
rect 583274 478046 583342 478102
rect 583398 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect -1916 477978 597980 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 6970 477978
rect 7026 477922 7094 477978
rect 7150 477922 7218 477978
rect 7274 477922 7342 477978
rect 7398 477922 24970 477978
rect 25026 477922 25094 477978
rect 25150 477922 25218 477978
rect 25274 477922 25342 477978
rect 25398 477922 42970 477978
rect 43026 477922 43094 477978
rect 43150 477922 43218 477978
rect 43274 477922 43342 477978
rect 43398 477922 60970 477978
rect 61026 477922 61094 477978
rect 61150 477922 61218 477978
rect 61274 477922 61342 477978
rect 61398 477922 69878 477978
rect 69934 477922 70002 477978
rect 70058 477922 78970 477978
rect 79026 477922 79094 477978
rect 79150 477922 79218 477978
rect 79274 477922 79342 477978
rect 79398 477922 96970 477978
rect 97026 477922 97094 477978
rect 97150 477922 97218 477978
rect 97274 477922 97342 477978
rect 97398 477922 100598 477978
rect 100654 477922 100722 477978
rect 100778 477922 131318 477978
rect 131374 477922 131442 477978
rect 131498 477922 162038 477978
rect 162094 477922 162162 477978
rect 162218 477922 192758 477978
rect 192814 477922 192882 477978
rect 192938 477922 223478 477978
rect 223534 477922 223602 477978
rect 223658 477922 254198 477978
rect 254254 477922 254322 477978
rect 254378 477922 284918 477978
rect 284974 477922 285042 477978
rect 285098 477922 315638 477978
rect 315694 477922 315762 477978
rect 315818 477922 346358 477978
rect 346414 477922 346482 477978
rect 346538 477922 377078 477978
rect 377134 477922 377202 477978
rect 377258 477922 407798 477978
rect 407854 477922 407922 477978
rect 407978 477922 438518 477978
rect 438574 477922 438642 477978
rect 438698 477922 469238 477978
rect 469294 477922 469362 477978
rect 469418 477922 499958 477978
rect 500014 477922 500082 477978
rect 500138 477922 530678 477978
rect 530734 477922 530802 477978
rect 530858 477922 564970 477978
rect 565026 477922 565094 477978
rect 565150 477922 565218 477978
rect 565274 477922 565342 477978
rect 565398 477922 582970 477978
rect 583026 477922 583094 477978
rect 583150 477922 583218 477978
rect 583274 477922 583342 477978
rect 583398 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect -1916 477826 597980 477922
rect -1916 472350 597980 472446
rect -1916 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 3250 472350
rect 3306 472294 3374 472350
rect 3430 472294 3498 472350
rect 3554 472294 3622 472350
rect 3678 472294 21250 472350
rect 21306 472294 21374 472350
rect 21430 472294 21498 472350
rect 21554 472294 21622 472350
rect 21678 472294 39250 472350
rect 39306 472294 39374 472350
rect 39430 472294 39498 472350
rect 39554 472294 39622 472350
rect 39678 472294 54518 472350
rect 54574 472294 54642 472350
rect 54698 472294 57250 472350
rect 57306 472294 57374 472350
rect 57430 472294 57498 472350
rect 57554 472294 57622 472350
rect 57678 472294 75250 472350
rect 75306 472294 75374 472350
rect 75430 472294 75498 472350
rect 75554 472294 75622 472350
rect 75678 472294 85238 472350
rect 85294 472294 85362 472350
rect 85418 472294 93250 472350
rect 93306 472294 93374 472350
rect 93430 472294 93498 472350
rect 93554 472294 93622 472350
rect 93678 472294 111250 472350
rect 111306 472294 111374 472350
rect 111430 472294 111498 472350
rect 111554 472294 111622 472350
rect 111678 472294 115958 472350
rect 116014 472294 116082 472350
rect 116138 472294 146678 472350
rect 146734 472294 146802 472350
rect 146858 472294 177398 472350
rect 177454 472294 177522 472350
rect 177578 472294 208118 472350
rect 208174 472294 208242 472350
rect 208298 472294 238838 472350
rect 238894 472294 238962 472350
rect 239018 472294 269558 472350
rect 269614 472294 269682 472350
rect 269738 472294 300278 472350
rect 300334 472294 300402 472350
rect 300458 472294 330998 472350
rect 331054 472294 331122 472350
rect 331178 472294 361718 472350
rect 361774 472294 361842 472350
rect 361898 472294 392438 472350
rect 392494 472294 392562 472350
rect 392618 472294 423158 472350
rect 423214 472294 423282 472350
rect 423338 472294 453878 472350
rect 453934 472294 454002 472350
rect 454058 472294 484598 472350
rect 484654 472294 484722 472350
rect 484778 472294 515318 472350
rect 515374 472294 515442 472350
rect 515498 472294 546038 472350
rect 546094 472294 546162 472350
rect 546218 472294 561250 472350
rect 561306 472294 561374 472350
rect 561430 472294 561498 472350
rect 561554 472294 561622 472350
rect 561678 472294 579250 472350
rect 579306 472294 579374 472350
rect 579430 472294 579498 472350
rect 579554 472294 579622 472350
rect 579678 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597980 472350
rect -1916 472226 597980 472294
rect -1916 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 3250 472226
rect 3306 472170 3374 472226
rect 3430 472170 3498 472226
rect 3554 472170 3622 472226
rect 3678 472170 21250 472226
rect 21306 472170 21374 472226
rect 21430 472170 21498 472226
rect 21554 472170 21622 472226
rect 21678 472170 39250 472226
rect 39306 472170 39374 472226
rect 39430 472170 39498 472226
rect 39554 472170 39622 472226
rect 39678 472170 54518 472226
rect 54574 472170 54642 472226
rect 54698 472170 57250 472226
rect 57306 472170 57374 472226
rect 57430 472170 57498 472226
rect 57554 472170 57622 472226
rect 57678 472170 75250 472226
rect 75306 472170 75374 472226
rect 75430 472170 75498 472226
rect 75554 472170 75622 472226
rect 75678 472170 85238 472226
rect 85294 472170 85362 472226
rect 85418 472170 93250 472226
rect 93306 472170 93374 472226
rect 93430 472170 93498 472226
rect 93554 472170 93622 472226
rect 93678 472170 111250 472226
rect 111306 472170 111374 472226
rect 111430 472170 111498 472226
rect 111554 472170 111622 472226
rect 111678 472170 115958 472226
rect 116014 472170 116082 472226
rect 116138 472170 146678 472226
rect 146734 472170 146802 472226
rect 146858 472170 177398 472226
rect 177454 472170 177522 472226
rect 177578 472170 208118 472226
rect 208174 472170 208242 472226
rect 208298 472170 238838 472226
rect 238894 472170 238962 472226
rect 239018 472170 269558 472226
rect 269614 472170 269682 472226
rect 269738 472170 300278 472226
rect 300334 472170 300402 472226
rect 300458 472170 330998 472226
rect 331054 472170 331122 472226
rect 331178 472170 361718 472226
rect 361774 472170 361842 472226
rect 361898 472170 392438 472226
rect 392494 472170 392562 472226
rect 392618 472170 423158 472226
rect 423214 472170 423282 472226
rect 423338 472170 453878 472226
rect 453934 472170 454002 472226
rect 454058 472170 484598 472226
rect 484654 472170 484722 472226
rect 484778 472170 515318 472226
rect 515374 472170 515442 472226
rect 515498 472170 546038 472226
rect 546094 472170 546162 472226
rect 546218 472170 561250 472226
rect 561306 472170 561374 472226
rect 561430 472170 561498 472226
rect 561554 472170 561622 472226
rect 561678 472170 579250 472226
rect 579306 472170 579374 472226
rect 579430 472170 579498 472226
rect 579554 472170 579622 472226
rect 579678 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597980 472226
rect -1916 472102 597980 472170
rect -1916 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 3250 472102
rect 3306 472046 3374 472102
rect 3430 472046 3498 472102
rect 3554 472046 3622 472102
rect 3678 472046 21250 472102
rect 21306 472046 21374 472102
rect 21430 472046 21498 472102
rect 21554 472046 21622 472102
rect 21678 472046 39250 472102
rect 39306 472046 39374 472102
rect 39430 472046 39498 472102
rect 39554 472046 39622 472102
rect 39678 472046 54518 472102
rect 54574 472046 54642 472102
rect 54698 472046 57250 472102
rect 57306 472046 57374 472102
rect 57430 472046 57498 472102
rect 57554 472046 57622 472102
rect 57678 472046 75250 472102
rect 75306 472046 75374 472102
rect 75430 472046 75498 472102
rect 75554 472046 75622 472102
rect 75678 472046 85238 472102
rect 85294 472046 85362 472102
rect 85418 472046 93250 472102
rect 93306 472046 93374 472102
rect 93430 472046 93498 472102
rect 93554 472046 93622 472102
rect 93678 472046 111250 472102
rect 111306 472046 111374 472102
rect 111430 472046 111498 472102
rect 111554 472046 111622 472102
rect 111678 472046 115958 472102
rect 116014 472046 116082 472102
rect 116138 472046 146678 472102
rect 146734 472046 146802 472102
rect 146858 472046 177398 472102
rect 177454 472046 177522 472102
rect 177578 472046 208118 472102
rect 208174 472046 208242 472102
rect 208298 472046 238838 472102
rect 238894 472046 238962 472102
rect 239018 472046 269558 472102
rect 269614 472046 269682 472102
rect 269738 472046 300278 472102
rect 300334 472046 300402 472102
rect 300458 472046 330998 472102
rect 331054 472046 331122 472102
rect 331178 472046 361718 472102
rect 361774 472046 361842 472102
rect 361898 472046 392438 472102
rect 392494 472046 392562 472102
rect 392618 472046 423158 472102
rect 423214 472046 423282 472102
rect 423338 472046 453878 472102
rect 453934 472046 454002 472102
rect 454058 472046 484598 472102
rect 484654 472046 484722 472102
rect 484778 472046 515318 472102
rect 515374 472046 515442 472102
rect 515498 472046 546038 472102
rect 546094 472046 546162 472102
rect 546218 472046 561250 472102
rect 561306 472046 561374 472102
rect 561430 472046 561498 472102
rect 561554 472046 561622 472102
rect 561678 472046 579250 472102
rect 579306 472046 579374 472102
rect 579430 472046 579498 472102
rect 579554 472046 579622 472102
rect 579678 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597980 472102
rect -1916 471978 597980 472046
rect -1916 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 3250 471978
rect 3306 471922 3374 471978
rect 3430 471922 3498 471978
rect 3554 471922 3622 471978
rect 3678 471922 21250 471978
rect 21306 471922 21374 471978
rect 21430 471922 21498 471978
rect 21554 471922 21622 471978
rect 21678 471922 39250 471978
rect 39306 471922 39374 471978
rect 39430 471922 39498 471978
rect 39554 471922 39622 471978
rect 39678 471922 54518 471978
rect 54574 471922 54642 471978
rect 54698 471922 57250 471978
rect 57306 471922 57374 471978
rect 57430 471922 57498 471978
rect 57554 471922 57622 471978
rect 57678 471922 75250 471978
rect 75306 471922 75374 471978
rect 75430 471922 75498 471978
rect 75554 471922 75622 471978
rect 75678 471922 85238 471978
rect 85294 471922 85362 471978
rect 85418 471922 93250 471978
rect 93306 471922 93374 471978
rect 93430 471922 93498 471978
rect 93554 471922 93622 471978
rect 93678 471922 111250 471978
rect 111306 471922 111374 471978
rect 111430 471922 111498 471978
rect 111554 471922 111622 471978
rect 111678 471922 115958 471978
rect 116014 471922 116082 471978
rect 116138 471922 146678 471978
rect 146734 471922 146802 471978
rect 146858 471922 177398 471978
rect 177454 471922 177522 471978
rect 177578 471922 208118 471978
rect 208174 471922 208242 471978
rect 208298 471922 238838 471978
rect 238894 471922 238962 471978
rect 239018 471922 269558 471978
rect 269614 471922 269682 471978
rect 269738 471922 300278 471978
rect 300334 471922 300402 471978
rect 300458 471922 330998 471978
rect 331054 471922 331122 471978
rect 331178 471922 361718 471978
rect 361774 471922 361842 471978
rect 361898 471922 392438 471978
rect 392494 471922 392562 471978
rect 392618 471922 423158 471978
rect 423214 471922 423282 471978
rect 423338 471922 453878 471978
rect 453934 471922 454002 471978
rect 454058 471922 484598 471978
rect 484654 471922 484722 471978
rect 484778 471922 515318 471978
rect 515374 471922 515442 471978
rect 515498 471922 546038 471978
rect 546094 471922 546162 471978
rect 546218 471922 561250 471978
rect 561306 471922 561374 471978
rect 561430 471922 561498 471978
rect 561554 471922 561622 471978
rect 561678 471922 579250 471978
rect 579306 471922 579374 471978
rect 579430 471922 579498 471978
rect 579554 471922 579622 471978
rect 579678 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597980 471978
rect -1916 471826 597980 471922
rect -1916 460350 597980 460446
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 6970 460350
rect 7026 460294 7094 460350
rect 7150 460294 7218 460350
rect 7274 460294 7342 460350
rect 7398 460294 24970 460350
rect 25026 460294 25094 460350
rect 25150 460294 25218 460350
rect 25274 460294 25342 460350
rect 25398 460294 42970 460350
rect 43026 460294 43094 460350
rect 43150 460294 43218 460350
rect 43274 460294 43342 460350
rect 43398 460294 60970 460350
rect 61026 460294 61094 460350
rect 61150 460294 61218 460350
rect 61274 460294 61342 460350
rect 61398 460294 69878 460350
rect 69934 460294 70002 460350
rect 70058 460294 78970 460350
rect 79026 460294 79094 460350
rect 79150 460294 79218 460350
rect 79274 460294 79342 460350
rect 79398 460294 96970 460350
rect 97026 460294 97094 460350
rect 97150 460294 97218 460350
rect 97274 460294 97342 460350
rect 97398 460294 100598 460350
rect 100654 460294 100722 460350
rect 100778 460294 131318 460350
rect 131374 460294 131442 460350
rect 131498 460294 162038 460350
rect 162094 460294 162162 460350
rect 162218 460294 192758 460350
rect 192814 460294 192882 460350
rect 192938 460294 223478 460350
rect 223534 460294 223602 460350
rect 223658 460294 254198 460350
rect 254254 460294 254322 460350
rect 254378 460294 284918 460350
rect 284974 460294 285042 460350
rect 285098 460294 315638 460350
rect 315694 460294 315762 460350
rect 315818 460294 346358 460350
rect 346414 460294 346482 460350
rect 346538 460294 377078 460350
rect 377134 460294 377202 460350
rect 377258 460294 407798 460350
rect 407854 460294 407922 460350
rect 407978 460294 438518 460350
rect 438574 460294 438642 460350
rect 438698 460294 469238 460350
rect 469294 460294 469362 460350
rect 469418 460294 499958 460350
rect 500014 460294 500082 460350
rect 500138 460294 530678 460350
rect 530734 460294 530802 460350
rect 530858 460294 564970 460350
rect 565026 460294 565094 460350
rect 565150 460294 565218 460350
rect 565274 460294 565342 460350
rect 565398 460294 582970 460350
rect 583026 460294 583094 460350
rect 583150 460294 583218 460350
rect 583274 460294 583342 460350
rect 583398 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect -1916 460226 597980 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 6970 460226
rect 7026 460170 7094 460226
rect 7150 460170 7218 460226
rect 7274 460170 7342 460226
rect 7398 460170 24970 460226
rect 25026 460170 25094 460226
rect 25150 460170 25218 460226
rect 25274 460170 25342 460226
rect 25398 460170 42970 460226
rect 43026 460170 43094 460226
rect 43150 460170 43218 460226
rect 43274 460170 43342 460226
rect 43398 460170 60970 460226
rect 61026 460170 61094 460226
rect 61150 460170 61218 460226
rect 61274 460170 61342 460226
rect 61398 460170 69878 460226
rect 69934 460170 70002 460226
rect 70058 460170 78970 460226
rect 79026 460170 79094 460226
rect 79150 460170 79218 460226
rect 79274 460170 79342 460226
rect 79398 460170 96970 460226
rect 97026 460170 97094 460226
rect 97150 460170 97218 460226
rect 97274 460170 97342 460226
rect 97398 460170 100598 460226
rect 100654 460170 100722 460226
rect 100778 460170 131318 460226
rect 131374 460170 131442 460226
rect 131498 460170 162038 460226
rect 162094 460170 162162 460226
rect 162218 460170 192758 460226
rect 192814 460170 192882 460226
rect 192938 460170 223478 460226
rect 223534 460170 223602 460226
rect 223658 460170 254198 460226
rect 254254 460170 254322 460226
rect 254378 460170 284918 460226
rect 284974 460170 285042 460226
rect 285098 460170 315638 460226
rect 315694 460170 315762 460226
rect 315818 460170 346358 460226
rect 346414 460170 346482 460226
rect 346538 460170 377078 460226
rect 377134 460170 377202 460226
rect 377258 460170 407798 460226
rect 407854 460170 407922 460226
rect 407978 460170 438518 460226
rect 438574 460170 438642 460226
rect 438698 460170 469238 460226
rect 469294 460170 469362 460226
rect 469418 460170 499958 460226
rect 500014 460170 500082 460226
rect 500138 460170 530678 460226
rect 530734 460170 530802 460226
rect 530858 460170 564970 460226
rect 565026 460170 565094 460226
rect 565150 460170 565218 460226
rect 565274 460170 565342 460226
rect 565398 460170 582970 460226
rect 583026 460170 583094 460226
rect 583150 460170 583218 460226
rect 583274 460170 583342 460226
rect 583398 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect -1916 460102 597980 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 6970 460102
rect 7026 460046 7094 460102
rect 7150 460046 7218 460102
rect 7274 460046 7342 460102
rect 7398 460046 24970 460102
rect 25026 460046 25094 460102
rect 25150 460046 25218 460102
rect 25274 460046 25342 460102
rect 25398 460046 42970 460102
rect 43026 460046 43094 460102
rect 43150 460046 43218 460102
rect 43274 460046 43342 460102
rect 43398 460046 60970 460102
rect 61026 460046 61094 460102
rect 61150 460046 61218 460102
rect 61274 460046 61342 460102
rect 61398 460046 69878 460102
rect 69934 460046 70002 460102
rect 70058 460046 78970 460102
rect 79026 460046 79094 460102
rect 79150 460046 79218 460102
rect 79274 460046 79342 460102
rect 79398 460046 96970 460102
rect 97026 460046 97094 460102
rect 97150 460046 97218 460102
rect 97274 460046 97342 460102
rect 97398 460046 100598 460102
rect 100654 460046 100722 460102
rect 100778 460046 131318 460102
rect 131374 460046 131442 460102
rect 131498 460046 162038 460102
rect 162094 460046 162162 460102
rect 162218 460046 192758 460102
rect 192814 460046 192882 460102
rect 192938 460046 223478 460102
rect 223534 460046 223602 460102
rect 223658 460046 254198 460102
rect 254254 460046 254322 460102
rect 254378 460046 284918 460102
rect 284974 460046 285042 460102
rect 285098 460046 315638 460102
rect 315694 460046 315762 460102
rect 315818 460046 346358 460102
rect 346414 460046 346482 460102
rect 346538 460046 377078 460102
rect 377134 460046 377202 460102
rect 377258 460046 407798 460102
rect 407854 460046 407922 460102
rect 407978 460046 438518 460102
rect 438574 460046 438642 460102
rect 438698 460046 469238 460102
rect 469294 460046 469362 460102
rect 469418 460046 499958 460102
rect 500014 460046 500082 460102
rect 500138 460046 530678 460102
rect 530734 460046 530802 460102
rect 530858 460046 564970 460102
rect 565026 460046 565094 460102
rect 565150 460046 565218 460102
rect 565274 460046 565342 460102
rect 565398 460046 582970 460102
rect 583026 460046 583094 460102
rect 583150 460046 583218 460102
rect 583274 460046 583342 460102
rect 583398 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect -1916 459978 597980 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 6970 459978
rect 7026 459922 7094 459978
rect 7150 459922 7218 459978
rect 7274 459922 7342 459978
rect 7398 459922 24970 459978
rect 25026 459922 25094 459978
rect 25150 459922 25218 459978
rect 25274 459922 25342 459978
rect 25398 459922 42970 459978
rect 43026 459922 43094 459978
rect 43150 459922 43218 459978
rect 43274 459922 43342 459978
rect 43398 459922 60970 459978
rect 61026 459922 61094 459978
rect 61150 459922 61218 459978
rect 61274 459922 61342 459978
rect 61398 459922 69878 459978
rect 69934 459922 70002 459978
rect 70058 459922 78970 459978
rect 79026 459922 79094 459978
rect 79150 459922 79218 459978
rect 79274 459922 79342 459978
rect 79398 459922 96970 459978
rect 97026 459922 97094 459978
rect 97150 459922 97218 459978
rect 97274 459922 97342 459978
rect 97398 459922 100598 459978
rect 100654 459922 100722 459978
rect 100778 459922 131318 459978
rect 131374 459922 131442 459978
rect 131498 459922 162038 459978
rect 162094 459922 162162 459978
rect 162218 459922 192758 459978
rect 192814 459922 192882 459978
rect 192938 459922 223478 459978
rect 223534 459922 223602 459978
rect 223658 459922 254198 459978
rect 254254 459922 254322 459978
rect 254378 459922 284918 459978
rect 284974 459922 285042 459978
rect 285098 459922 315638 459978
rect 315694 459922 315762 459978
rect 315818 459922 346358 459978
rect 346414 459922 346482 459978
rect 346538 459922 377078 459978
rect 377134 459922 377202 459978
rect 377258 459922 407798 459978
rect 407854 459922 407922 459978
rect 407978 459922 438518 459978
rect 438574 459922 438642 459978
rect 438698 459922 469238 459978
rect 469294 459922 469362 459978
rect 469418 459922 499958 459978
rect 500014 459922 500082 459978
rect 500138 459922 530678 459978
rect 530734 459922 530802 459978
rect 530858 459922 564970 459978
rect 565026 459922 565094 459978
rect 565150 459922 565218 459978
rect 565274 459922 565342 459978
rect 565398 459922 582970 459978
rect 583026 459922 583094 459978
rect 583150 459922 583218 459978
rect 583274 459922 583342 459978
rect 583398 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect -1916 459826 597980 459922
rect -1916 454350 597980 454446
rect -1916 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 3250 454350
rect 3306 454294 3374 454350
rect 3430 454294 3498 454350
rect 3554 454294 3622 454350
rect 3678 454294 21250 454350
rect 21306 454294 21374 454350
rect 21430 454294 21498 454350
rect 21554 454294 21622 454350
rect 21678 454294 39250 454350
rect 39306 454294 39374 454350
rect 39430 454294 39498 454350
rect 39554 454294 39622 454350
rect 39678 454294 54518 454350
rect 54574 454294 54642 454350
rect 54698 454294 57250 454350
rect 57306 454294 57374 454350
rect 57430 454294 57498 454350
rect 57554 454294 57622 454350
rect 57678 454294 75250 454350
rect 75306 454294 75374 454350
rect 75430 454294 75498 454350
rect 75554 454294 75622 454350
rect 75678 454294 85238 454350
rect 85294 454294 85362 454350
rect 85418 454294 93250 454350
rect 93306 454294 93374 454350
rect 93430 454294 93498 454350
rect 93554 454294 93622 454350
rect 93678 454294 111250 454350
rect 111306 454294 111374 454350
rect 111430 454294 111498 454350
rect 111554 454294 111622 454350
rect 111678 454294 115958 454350
rect 116014 454294 116082 454350
rect 116138 454294 146678 454350
rect 146734 454294 146802 454350
rect 146858 454294 177398 454350
rect 177454 454294 177522 454350
rect 177578 454294 208118 454350
rect 208174 454294 208242 454350
rect 208298 454294 238838 454350
rect 238894 454294 238962 454350
rect 239018 454294 269558 454350
rect 269614 454294 269682 454350
rect 269738 454294 300278 454350
rect 300334 454294 300402 454350
rect 300458 454294 330998 454350
rect 331054 454294 331122 454350
rect 331178 454294 361718 454350
rect 361774 454294 361842 454350
rect 361898 454294 392438 454350
rect 392494 454294 392562 454350
rect 392618 454294 423158 454350
rect 423214 454294 423282 454350
rect 423338 454294 453878 454350
rect 453934 454294 454002 454350
rect 454058 454294 484598 454350
rect 484654 454294 484722 454350
rect 484778 454294 515318 454350
rect 515374 454294 515442 454350
rect 515498 454294 546038 454350
rect 546094 454294 546162 454350
rect 546218 454294 561250 454350
rect 561306 454294 561374 454350
rect 561430 454294 561498 454350
rect 561554 454294 561622 454350
rect 561678 454294 579250 454350
rect 579306 454294 579374 454350
rect 579430 454294 579498 454350
rect 579554 454294 579622 454350
rect 579678 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597980 454350
rect -1916 454226 597980 454294
rect -1916 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 3250 454226
rect 3306 454170 3374 454226
rect 3430 454170 3498 454226
rect 3554 454170 3622 454226
rect 3678 454170 21250 454226
rect 21306 454170 21374 454226
rect 21430 454170 21498 454226
rect 21554 454170 21622 454226
rect 21678 454170 39250 454226
rect 39306 454170 39374 454226
rect 39430 454170 39498 454226
rect 39554 454170 39622 454226
rect 39678 454170 54518 454226
rect 54574 454170 54642 454226
rect 54698 454170 57250 454226
rect 57306 454170 57374 454226
rect 57430 454170 57498 454226
rect 57554 454170 57622 454226
rect 57678 454170 75250 454226
rect 75306 454170 75374 454226
rect 75430 454170 75498 454226
rect 75554 454170 75622 454226
rect 75678 454170 85238 454226
rect 85294 454170 85362 454226
rect 85418 454170 93250 454226
rect 93306 454170 93374 454226
rect 93430 454170 93498 454226
rect 93554 454170 93622 454226
rect 93678 454170 111250 454226
rect 111306 454170 111374 454226
rect 111430 454170 111498 454226
rect 111554 454170 111622 454226
rect 111678 454170 115958 454226
rect 116014 454170 116082 454226
rect 116138 454170 146678 454226
rect 146734 454170 146802 454226
rect 146858 454170 177398 454226
rect 177454 454170 177522 454226
rect 177578 454170 208118 454226
rect 208174 454170 208242 454226
rect 208298 454170 238838 454226
rect 238894 454170 238962 454226
rect 239018 454170 269558 454226
rect 269614 454170 269682 454226
rect 269738 454170 300278 454226
rect 300334 454170 300402 454226
rect 300458 454170 330998 454226
rect 331054 454170 331122 454226
rect 331178 454170 361718 454226
rect 361774 454170 361842 454226
rect 361898 454170 392438 454226
rect 392494 454170 392562 454226
rect 392618 454170 423158 454226
rect 423214 454170 423282 454226
rect 423338 454170 453878 454226
rect 453934 454170 454002 454226
rect 454058 454170 484598 454226
rect 484654 454170 484722 454226
rect 484778 454170 515318 454226
rect 515374 454170 515442 454226
rect 515498 454170 546038 454226
rect 546094 454170 546162 454226
rect 546218 454170 561250 454226
rect 561306 454170 561374 454226
rect 561430 454170 561498 454226
rect 561554 454170 561622 454226
rect 561678 454170 579250 454226
rect 579306 454170 579374 454226
rect 579430 454170 579498 454226
rect 579554 454170 579622 454226
rect 579678 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597980 454226
rect -1916 454102 597980 454170
rect -1916 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 3250 454102
rect 3306 454046 3374 454102
rect 3430 454046 3498 454102
rect 3554 454046 3622 454102
rect 3678 454046 21250 454102
rect 21306 454046 21374 454102
rect 21430 454046 21498 454102
rect 21554 454046 21622 454102
rect 21678 454046 39250 454102
rect 39306 454046 39374 454102
rect 39430 454046 39498 454102
rect 39554 454046 39622 454102
rect 39678 454046 54518 454102
rect 54574 454046 54642 454102
rect 54698 454046 57250 454102
rect 57306 454046 57374 454102
rect 57430 454046 57498 454102
rect 57554 454046 57622 454102
rect 57678 454046 75250 454102
rect 75306 454046 75374 454102
rect 75430 454046 75498 454102
rect 75554 454046 75622 454102
rect 75678 454046 85238 454102
rect 85294 454046 85362 454102
rect 85418 454046 93250 454102
rect 93306 454046 93374 454102
rect 93430 454046 93498 454102
rect 93554 454046 93622 454102
rect 93678 454046 111250 454102
rect 111306 454046 111374 454102
rect 111430 454046 111498 454102
rect 111554 454046 111622 454102
rect 111678 454046 115958 454102
rect 116014 454046 116082 454102
rect 116138 454046 146678 454102
rect 146734 454046 146802 454102
rect 146858 454046 177398 454102
rect 177454 454046 177522 454102
rect 177578 454046 208118 454102
rect 208174 454046 208242 454102
rect 208298 454046 238838 454102
rect 238894 454046 238962 454102
rect 239018 454046 269558 454102
rect 269614 454046 269682 454102
rect 269738 454046 300278 454102
rect 300334 454046 300402 454102
rect 300458 454046 330998 454102
rect 331054 454046 331122 454102
rect 331178 454046 361718 454102
rect 361774 454046 361842 454102
rect 361898 454046 392438 454102
rect 392494 454046 392562 454102
rect 392618 454046 423158 454102
rect 423214 454046 423282 454102
rect 423338 454046 453878 454102
rect 453934 454046 454002 454102
rect 454058 454046 484598 454102
rect 484654 454046 484722 454102
rect 484778 454046 515318 454102
rect 515374 454046 515442 454102
rect 515498 454046 546038 454102
rect 546094 454046 546162 454102
rect 546218 454046 561250 454102
rect 561306 454046 561374 454102
rect 561430 454046 561498 454102
rect 561554 454046 561622 454102
rect 561678 454046 579250 454102
rect 579306 454046 579374 454102
rect 579430 454046 579498 454102
rect 579554 454046 579622 454102
rect 579678 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597980 454102
rect -1916 453978 597980 454046
rect -1916 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 3250 453978
rect 3306 453922 3374 453978
rect 3430 453922 3498 453978
rect 3554 453922 3622 453978
rect 3678 453922 21250 453978
rect 21306 453922 21374 453978
rect 21430 453922 21498 453978
rect 21554 453922 21622 453978
rect 21678 453922 39250 453978
rect 39306 453922 39374 453978
rect 39430 453922 39498 453978
rect 39554 453922 39622 453978
rect 39678 453922 54518 453978
rect 54574 453922 54642 453978
rect 54698 453922 57250 453978
rect 57306 453922 57374 453978
rect 57430 453922 57498 453978
rect 57554 453922 57622 453978
rect 57678 453922 75250 453978
rect 75306 453922 75374 453978
rect 75430 453922 75498 453978
rect 75554 453922 75622 453978
rect 75678 453922 85238 453978
rect 85294 453922 85362 453978
rect 85418 453922 93250 453978
rect 93306 453922 93374 453978
rect 93430 453922 93498 453978
rect 93554 453922 93622 453978
rect 93678 453922 111250 453978
rect 111306 453922 111374 453978
rect 111430 453922 111498 453978
rect 111554 453922 111622 453978
rect 111678 453922 115958 453978
rect 116014 453922 116082 453978
rect 116138 453922 146678 453978
rect 146734 453922 146802 453978
rect 146858 453922 177398 453978
rect 177454 453922 177522 453978
rect 177578 453922 208118 453978
rect 208174 453922 208242 453978
rect 208298 453922 238838 453978
rect 238894 453922 238962 453978
rect 239018 453922 269558 453978
rect 269614 453922 269682 453978
rect 269738 453922 300278 453978
rect 300334 453922 300402 453978
rect 300458 453922 330998 453978
rect 331054 453922 331122 453978
rect 331178 453922 361718 453978
rect 361774 453922 361842 453978
rect 361898 453922 392438 453978
rect 392494 453922 392562 453978
rect 392618 453922 423158 453978
rect 423214 453922 423282 453978
rect 423338 453922 453878 453978
rect 453934 453922 454002 453978
rect 454058 453922 484598 453978
rect 484654 453922 484722 453978
rect 484778 453922 515318 453978
rect 515374 453922 515442 453978
rect 515498 453922 546038 453978
rect 546094 453922 546162 453978
rect 546218 453922 561250 453978
rect 561306 453922 561374 453978
rect 561430 453922 561498 453978
rect 561554 453922 561622 453978
rect 561678 453922 579250 453978
rect 579306 453922 579374 453978
rect 579430 453922 579498 453978
rect 579554 453922 579622 453978
rect 579678 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597980 453978
rect -1916 453826 597980 453922
rect -1916 442350 597980 442446
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 6970 442350
rect 7026 442294 7094 442350
rect 7150 442294 7218 442350
rect 7274 442294 7342 442350
rect 7398 442294 24970 442350
rect 25026 442294 25094 442350
rect 25150 442294 25218 442350
rect 25274 442294 25342 442350
rect 25398 442294 42970 442350
rect 43026 442294 43094 442350
rect 43150 442294 43218 442350
rect 43274 442294 43342 442350
rect 43398 442294 60970 442350
rect 61026 442294 61094 442350
rect 61150 442294 61218 442350
rect 61274 442294 61342 442350
rect 61398 442294 69878 442350
rect 69934 442294 70002 442350
rect 70058 442294 78970 442350
rect 79026 442294 79094 442350
rect 79150 442294 79218 442350
rect 79274 442294 79342 442350
rect 79398 442294 96970 442350
rect 97026 442294 97094 442350
rect 97150 442294 97218 442350
rect 97274 442294 97342 442350
rect 97398 442294 100598 442350
rect 100654 442294 100722 442350
rect 100778 442294 131318 442350
rect 131374 442294 131442 442350
rect 131498 442294 162038 442350
rect 162094 442294 162162 442350
rect 162218 442294 192758 442350
rect 192814 442294 192882 442350
rect 192938 442294 223478 442350
rect 223534 442294 223602 442350
rect 223658 442294 254198 442350
rect 254254 442294 254322 442350
rect 254378 442294 284918 442350
rect 284974 442294 285042 442350
rect 285098 442294 315638 442350
rect 315694 442294 315762 442350
rect 315818 442294 346358 442350
rect 346414 442294 346482 442350
rect 346538 442294 377078 442350
rect 377134 442294 377202 442350
rect 377258 442294 407798 442350
rect 407854 442294 407922 442350
rect 407978 442294 438518 442350
rect 438574 442294 438642 442350
rect 438698 442294 469238 442350
rect 469294 442294 469362 442350
rect 469418 442294 499958 442350
rect 500014 442294 500082 442350
rect 500138 442294 530678 442350
rect 530734 442294 530802 442350
rect 530858 442294 564970 442350
rect 565026 442294 565094 442350
rect 565150 442294 565218 442350
rect 565274 442294 565342 442350
rect 565398 442294 582970 442350
rect 583026 442294 583094 442350
rect 583150 442294 583218 442350
rect 583274 442294 583342 442350
rect 583398 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect -1916 442226 597980 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 6970 442226
rect 7026 442170 7094 442226
rect 7150 442170 7218 442226
rect 7274 442170 7342 442226
rect 7398 442170 24970 442226
rect 25026 442170 25094 442226
rect 25150 442170 25218 442226
rect 25274 442170 25342 442226
rect 25398 442170 42970 442226
rect 43026 442170 43094 442226
rect 43150 442170 43218 442226
rect 43274 442170 43342 442226
rect 43398 442170 60970 442226
rect 61026 442170 61094 442226
rect 61150 442170 61218 442226
rect 61274 442170 61342 442226
rect 61398 442170 69878 442226
rect 69934 442170 70002 442226
rect 70058 442170 78970 442226
rect 79026 442170 79094 442226
rect 79150 442170 79218 442226
rect 79274 442170 79342 442226
rect 79398 442170 96970 442226
rect 97026 442170 97094 442226
rect 97150 442170 97218 442226
rect 97274 442170 97342 442226
rect 97398 442170 100598 442226
rect 100654 442170 100722 442226
rect 100778 442170 131318 442226
rect 131374 442170 131442 442226
rect 131498 442170 162038 442226
rect 162094 442170 162162 442226
rect 162218 442170 192758 442226
rect 192814 442170 192882 442226
rect 192938 442170 223478 442226
rect 223534 442170 223602 442226
rect 223658 442170 254198 442226
rect 254254 442170 254322 442226
rect 254378 442170 284918 442226
rect 284974 442170 285042 442226
rect 285098 442170 315638 442226
rect 315694 442170 315762 442226
rect 315818 442170 346358 442226
rect 346414 442170 346482 442226
rect 346538 442170 377078 442226
rect 377134 442170 377202 442226
rect 377258 442170 407798 442226
rect 407854 442170 407922 442226
rect 407978 442170 438518 442226
rect 438574 442170 438642 442226
rect 438698 442170 469238 442226
rect 469294 442170 469362 442226
rect 469418 442170 499958 442226
rect 500014 442170 500082 442226
rect 500138 442170 530678 442226
rect 530734 442170 530802 442226
rect 530858 442170 564970 442226
rect 565026 442170 565094 442226
rect 565150 442170 565218 442226
rect 565274 442170 565342 442226
rect 565398 442170 582970 442226
rect 583026 442170 583094 442226
rect 583150 442170 583218 442226
rect 583274 442170 583342 442226
rect 583398 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect -1916 442102 597980 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 6970 442102
rect 7026 442046 7094 442102
rect 7150 442046 7218 442102
rect 7274 442046 7342 442102
rect 7398 442046 24970 442102
rect 25026 442046 25094 442102
rect 25150 442046 25218 442102
rect 25274 442046 25342 442102
rect 25398 442046 42970 442102
rect 43026 442046 43094 442102
rect 43150 442046 43218 442102
rect 43274 442046 43342 442102
rect 43398 442046 60970 442102
rect 61026 442046 61094 442102
rect 61150 442046 61218 442102
rect 61274 442046 61342 442102
rect 61398 442046 69878 442102
rect 69934 442046 70002 442102
rect 70058 442046 78970 442102
rect 79026 442046 79094 442102
rect 79150 442046 79218 442102
rect 79274 442046 79342 442102
rect 79398 442046 96970 442102
rect 97026 442046 97094 442102
rect 97150 442046 97218 442102
rect 97274 442046 97342 442102
rect 97398 442046 100598 442102
rect 100654 442046 100722 442102
rect 100778 442046 131318 442102
rect 131374 442046 131442 442102
rect 131498 442046 162038 442102
rect 162094 442046 162162 442102
rect 162218 442046 192758 442102
rect 192814 442046 192882 442102
rect 192938 442046 223478 442102
rect 223534 442046 223602 442102
rect 223658 442046 254198 442102
rect 254254 442046 254322 442102
rect 254378 442046 284918 442102
rect 284974 442046 285042 442102
rect 285098 442046 315638 442102
rect 315694 442046 315762 442102
rect 315818 442046 346358 442102
rect 346414 442046 346482 442102
rect 346538 442046 377078 442102
rect 377134 442046 377202 442102
rect 377258 442046 407798 442102
rect 407854 442046 407922 442102
rect 407978 442046 438518 442102
rect 438574 442046 438642 442102
rect 438698 442046 469238 442102
rect 469294 442046 469362 442102
rect 469418 442046 499958 442102
rect 500014 442046 500082 442102
rect 500138 442046 530678 442102
rect 530734 442046 530802 442102
rect 530858 442046 564970 442102
rect 565026 442046 565094 442102
rect 565150 442046 565218 442102
rect 565274 442046 565342 442102
rect 565398 442046 582970 442102
rect 583026 442046 583094 442102
rect 583150 442046 583218 442102
rect 583274 442046 583342 442102
rect 583398 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect -1916 441978 597980 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 6970 441978
rect 7026 441922 7094 441978
rect 7150 441922 7218 441978
rect 7274 441922 7342 441978
rect 7398 441922 24970 441978
rect 25026 441922 25094 441978
rect 25150 441922 25218 441978
rect 25274 441922 25342 441978
rect 25398 441922 42970 441978
rect 43026 441922 43094 441978
rect 43150 441922 43218 441978
rect 43274 441922 43342 441978
rect 43398 441922 60970 441978
rect 61026 441922 61094 441978
rect 61150 441922 61218 441978
rect 61274 441922 61342 441978
rect 61398 441922 69878 441978
rect 69934 441922 70002 441978
rect 70058 441922 78970 441978
rect 79026 441922 79094 441978
rect 79150 441922 79218 441978
rect 79274 441922 79342 441978
rect 79398 441922 96970 441978
rect 97026 441922 97094 441978
rect 97150 441922 97218 441978
rect 97274 441922 97342 441978
rect 97398 441922 100598 441978
rect 100654 441922 100722 441978
rect 100778 441922 131318 441978
rect 131374 441922 131442 441978
rect 131498 441922 162038 441978
rect 162094 441922 162162 441978
rect 162218 441922 192758 441978
rect 192814 441922 192882 441978
rect 192938 441922 223478 441978
rect 223534 441922 223602 441978
rect 223658 441922 254198 441978
rect 254254 441922 254322 441978
rect 254378 441922 284918 441978
rect 284974 441922 285042 441978
rect 285098 441922 315638 441978
rect 315694 441922 315762 441978
rect 315818 441922 346358 441978
rect 346414 441922 346482 441978
rect 346538 441922 377078 441978
rect 377134 441922 377202 441978
rect 377258 441922 407798 441978
rect 407854 441922 407922 441978
rect 407978 441922 438518 441978
rect 438574 441922 438642 441978
rect 438698 441922 469238 441978
rect 469294 441922 469362 441978
rect 469418 441922 499958 441978
rect 500014 441922 500082 441978
rect 500138 441922 530678 441978
rect 530734 441922 530802 441978
rect 530858 441922 564970 441978
rect 565026 441922 565094 441978
rect 565150 441922 565218 441978
rect 565274 441922 565342 441978
rect 565398 441922 582970 441978
rect 583026 441922 583094 441978
rect 583150 441922 583218 441978
rect 583274 441922 583342 441978
rect 583398 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect -1916 441826 597980 441922
rect -1916 436350 597980 436446
rect -1916 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 3250 436350
rect 3306 436294 3374 436350
rect 3430 436294 3498 436350
rect 3554 436294 3622 436350
rect 3678 436294 21250 436350
rect 21306 436294 21374 436350
rect 21430 436294 21498 436350
rect 21554 436294 21622 436350
rect 21678 436294 39250 436350
rect 39306 436294 39374 436350
rect 39430 436294 39498 436350
rect 39554 436294 39622 436350
rect 39678 436294 54518 436350
rect 54574 436294 54642 436350
rect 54698 436294 57250 436350
rect 57306 436294 57374 436350
rect 57430 436294 57498 436350
rect 57554 436294 57622 436350
rect 57678 436294 75250 436350
rect 75306 436294 75374 436350
rect 75430 436294 75498 436350
rect 75554 436294 75622 436350
rect 75678 436294 85238 436350
rect 85294 436294 85362 436350
rect 85418 436294 93250 436350
rect 93306 436294 93374 436350
rect 93430 436294 93498 436350
rect 93554 436294 93622 436350
rect 93678 436294 111250 436350
rect 111306 436294 111374 436350
rect 111430 436294 111498 436350
rect 111554 436294 111622 436350
rect 111678 436294 115958 436350
rect 116014 436294 116082 436350
rect 116138 436294 146678 436350
rect 146734 436294 146802 436350
rect 146858 436294 177398 436350
rect 177454 436294 177522 436350
rect 177578 436294 208118 436350
rect 208174 436294 208242 436350
rect 208298 436294 238838 436350
rect 238894 436294 238962 436350
rect 239018 436294 269558 436350
rect 269614 436294 269682 436350
rect 269738 436294 300278 436350
rect 300334 436294 300402 436350
rect 300458 436294 330998 436350
rect 331054 436294 331122 436350
rect 331178 436294 361718 436350
rect 361774 436294 361842 436350
rect 361898 436294 392438 436350
rect 392494 436294 392562 436350
rect 392618 436294 423158 436350
rect 423214 436294 423282 436350
rect 423338 436294 453878 436350
rect 453934 436294 454002 436350
rect 454058 436294 484598 436350
rect 484654 436294 484722 436350
rect 484778 436294 515318 436350
rect 515374 436294 515442 436350
rect 515498 436294 546038 436350
rect 546094 436294 546162 436350
rect 546218 436294 561250 436350
rect 561306 436294 561374 436350
rect 561430 436294 561498 436350
rect 561554 436294 561622 436350
rect 561678 436294 579250 436350
rect 579306 436294 579374 436350
rect 579430 436294 579498 436350
rect 579554 436294 579622 436350
rect 579678 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597980 436350
rect -1916 436226 597980 436294
rect -1916 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 3250 436226
rect 3306 436170 3374 436226
rect 3430 436170 3498 436226
rect 3554 436170 3622 436226
rect 3678 436170 21250 436226
rect 21306 436170 21374 436226
rect 21430 436170 21498 436226
rect 21554 436170 21622 436226
rect 21678 436170 39250 436226
rect 39306 436170 39374 436226
rect 39430 436170 39498 436226
rect 39554 436170 39622 436226
rect 39678 436170 54518 436226
rect 54574 436170 54642 436226
rect 54698 436170 57250 436226
rect 57306 436170 57374 436226
rect 57430 436170 57498 436226
rect 57554 436170 57622 436226
rect 57678 436170 75250 436226
rect 75306 436170 75374 436226
rect 75430 436170 75498 436226
rect 75554 436170 75622 436226
rect 75678 436170 85238 436226
rect 85294 436170 85362 436226
rect 85418 436170 93250 436226
rect 93306 436170 93374 436226
rect 93430 436170 93498 436226
rect 93554 436170 93622 436226
rect 93678 436170 111250 436226
rect 111306 436170 111374 436226
rect 111430 436170 111498 436226
rect 111554 436170 111622 436226
rect 111678 436170 115958 436226
rect 116014 436170 116082 436226
rect 116138 436170 146678 436226
rect 146734 436170 146802 436226
rect 146858 436170 177398 436226
rect 177454 436170 177522 436226
rect 177578 436170 208118 436226
rect 208174 436170 208242 436226
rect 208298 436170 238838 436226
rect 238894 436170 238962 436226
rect 239018 436170 269558 436226
rect 269614 436170 269682 436226
rect 269738 436170 300278 436226
rect 300334 436170 300402 436226
rect 300458 436170 330998 436226
rect 331054 436170 331122 436226
rect 331178 436170 361718 436226
rect 361774 436170 361842 436226
rect 361898 436170 392438 436226
rect 392494 436170 392562 436226
rect 392618 436170 423158 436226
rect 423214 436170 423282 436226
rect 423338 436170 453878 436226
rect 453934 436170 454002 436226
rect 454058 436170 484598 436226
rect 484654 436170 484722 436226
rect 484778 436170 515318 436226
rect 515374 436170 515442 436226
rect 515498 436170 546038 436226
rect 546094 436170 546162 436226
rect 546218 436170 561250 436226
rect 561306 436170 561374 436226
rect 561430 436170 561498 436226
rect 561554 436170 561622 436226
rect 561678 436170 579250 436226
rect 579306 436170 579374 436226
rect 579430 436170 579498 436226
rect 579554 436170 579622 436226
rect 579678 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597980 436226
rect -1916 436102 597980 436170
rect -1916 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 3250 436102
rect 3306 436046 3374 436102
rect 3430 436046 3498 436102
rect 3554 436046 3622 436102
rect 3678 436046 21250 436102
rect 21306 436046 21374 436102
rect 21430 436046 21498 436102
rect 21554 436046 21622 436102
rect 21678 436046 39250 436102
rect 39306 436046 39374 436102
rect 39430 436046 39498 436102
rect 39554 436046 39622 436102
rect 39678 436046 54518 436102
rect 54574 436046 54642 436102
rect 54698 436046 57250 436102
rect 57306 436046 57374 436102
rect 57430 436046 57498 436102
rect 57554 436046 57622 436102
rect 57678 436046 75250 436102
rect 75306 436046 75374 436102
rect 75430 436046 75498 436102
rect 75554 436046 75622 436102
rect 75678 436046 85238 436102
rect 85294 436046 85362 436102
rect 85418 436046 93250 436102
rect 93306 436046 93374 436102
rect 93430 436046 93498 436102
rect 93554 436046 93622 436102
rect 93678 436046 111250 436102
rect 111306 436046 111374 436102
rect 111430 436046 111498 436102
rect 111554 436046 111622 436102
rect 111678 436046 115958 436102
rect 116014 436046 116082 436102
rect 116138 436046 146678 436102
rect 146734 436046 146802 436102
rect 146858 436046 177398 436102
rect 177454 436046 177522 436102
rect 177578 436046 208118 436102
rect 208174 436046 208242 436102
rect 208298 436046 238838 436102
rect 238894 436046 238962 436102
rect 239018 436046 269558 436102
rect 269614 436046 269682 436102
rect 269738 436046 300278 436102
rect 300334 436046 300402 436102
rect 300458 436046 330998 436102
rect 331054 436046 331122 436102
rect 331178 436046 361718 436102
rect 361774 436046 361842 436102
rect 361898 436046 392438 436102
rect 392494 436046 392562 436102
rect 392618 436046 423158 436102
rect 423214 436046 423282 436102
rect 423338 436046 453878 436102
rect 453934 436046 454002 436102
rect 454058 436046 484598 436102
rect 484654 436046 484722 436102
rect 484778 436046 515318 436102
rect 515374 436046 515442 436102
rect 515498 436046 546038 436102
rect 546094 436046 546162 436102
rect 546218 436046 561250 436102
rect 561306 436046 561374 436102
rect 561430 436046 561498 436102
rect 561554 436046 561622 436102
rect 561678 436046 579250 436102
rect 579306 436046 579374 436102
rect 579430 436046 579498 436102
rect 579554 436046 579622 436102
rect 579678 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597980 436102
rect -1916 435978 597980 436046
rect -1916 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 3250 435978
rect 3306 435922 3374 435978
rect 3430 435922 3498 435978
rect 3554 435922 3622 435978
rect 3678 435922 21250 435978
rect 21306 435922 21374 435978
rect 21430 435922 21498 435978
rect 21554 435922 21622 435978
rect 21678 435922 39250 435978
rect 39306 435922 39374 435978
rect 39430 435922 39498 435978
rect 39554 435922 39622 435978
rect 39678 435922 54518 435978
rect 54574 435922 54642 435978
rect 54698 435922 57250 435978
rect 57306 435922 57374 435978
rect 57430 435922 57498 435978
rect 57554 435922 57622 435978
rect 57678 435922 75250 435978
rect 75306 435922 75374 435978
rect 75430 435922 75498 435978
rect 75554 435922 75622 435978
rect 75678 435922 85238 435978
rect 85294 435922 85362 435978
rect 85418 435922 93250 435978
rect 93306 435922 93374 435978
rect 93430 435922 93498 435978
rect 93554 435922 93622 435978
rect 93678 435922 111250 435978
rect 111306 435922 111374 435978
rect 111430 435922 111498 435978
rect 111554 435922 111622 435978
rect 111678 435922 115958 435978
rect 116014 435922 116082 435978
rect 116138 435922 146678 435978
rect 146734 435922 146802 435978
rect 146858 435922 177398 435978
rect 177454 435922 177522 435978
rect 177578 435922 208118 435978
rect 208174 435922 208242 435978
rect 208298 435922 238838 435978
rect 238894 435922 238962 435978
rect 239018 435922 269558 435978
rect 269614 435922 269682 435978
rect 269738 435922 300278 435978
rect 300334 435922 300402 435978
rect 300458 435922 330998 435978
rect 331054 435922 331122 435978
rect 331178 435922 361718 435978
rect 361774 435922 361842 435978
rect 361898 435922 392438 435978
rect 392494 435922 392562 435978
rect 392618 435922 423158 435978
rect 423214 435922 423282 435978
rect 423338 435922 453878 435978
rect 453934 435922 454002 435978
rect 454058 435922 484598 435978
rect 484654 435922 484722 435978
rect 484778 435922 515318 435978
rect 515374 435922 515442 435978
rect 515498 435922 546038 435978
rect 546094 435922 546162 435978
rect 546218 435922 561250 435978
rect 561306 435922 561374 435978
rect 561430 435922 561498 435978
rect 561554 435922 561622 435978
rect 561678 435922 579250 435978
rect 579306 435922 579374 435978
rect 579430 435922 579498 435978
rect 579554 435922 579622 435978
rect 579678 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597980 435978
rect -1916 435826 597980 435922
rect -1916 424350 597980 424446
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 6970 424350
rect 7026 424294 7094 424350
rect 7150 424294 7218 424350
rect 7274 424294 7342 424350
rect 7398 424294 24970 424350
rect 25026 424294 25094 424350
rect 25150 424294 25218 424350
rect 25274 424294 25342 424350
rect 25398 424294 42970 424350
rect 43026 424294 43094 424350
rect 43150 424294 43218 424350
rect 43274 424294 43342 424350
rect 43398 424294 60970 424350
rect 61026 424294 61094 424350
rect 61150 424294 61218 424350
rect 61274 424294 61342 424350
rect 61398 424294 69878 424350
rect 69934 424294 70002 424350
rect 70058 424294 78970 424350
rect 79026 424294 79094 424350
rect 79150 424294 79218 424350
rect 79274 424294 79342 424350
rect 79398 424294 96970 424350
rect 97026 424294 97094 424350
rect 97150 424294 97218 424350
rect 97274 424294 97342 424350
rect 97398 424294 100598 424350
rect 100654 424294 100722 424350
rect 100778 424294 131318 424350
rect 131374 424294 131442 424350
rect 131498 424294 162038 424350
rect 162094 424294 162162 424350
rect 162218 424294 192758 424350
rect 192814 424294 192882 424350
rect 192938 424294 223478 424350
rect 223534 424294 223602 424350
rect 223658 424294 254198 424350
rect 254254 424294 254322 424350
rect 254378 424294 284918 424350
rect 284974 424294 285042 424350
rect 285098 424294 315638 424350
rect 315694 424294 315762 424350
rect 315818 424294 346358 424350
rect 346414 424294 346482 424350
rect 346538 424294 377078 424350
rect 377134 424294 377202 424350
rect 377258 424294 407798 424350
rect 407854 424294 407922 424350
rect 407978 424294 438518 424350
rect 438574 424294 438642 424350
rect 438698 424294 469238 424350
rect 469294 424294 469362 424350
rect 469418 424294 499958 424350
rect 500014 424294 500082 424350
rect 500138 424294 530678 424350
rect 530734 424294 530802 424350
rect 530858 424294 564970 424350
rect 565026 424294 565094 424350
rect 565150 424294 565218 424350
rect 565274 424294 565342 424350
rect 565398 424294 582970 424350
rect 583026 424294 583094 424350
rect 583150 424294 583218 424350
rect 583274 424294 583342 424350
rect 583398 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect -1916 424226 597980 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 6970 424226
rect 7026 424170 7094 424226
rect 7150 424170 7218 424226
rect 7274 424170 7342 424226
rect 7398 424170 24970 424226
rect 25026 424170 25094 424226
rect 25150 424170 25218 424226
rect 25274 424170 25342 424226
rect 25398 424170 42970 424226
rect 43026 424170 43094 424226
rect 43150 424170 43218 424226
rect 43274 424170 43342 424226
rect 43398 424170 60970 424226
rect 61026 424170 61094 424226
rect 61150 424170 61218 424226
rect 61274 424170 61342 424226
rect 61398 424170 69878 424226
rect 69934 424170 70002 424226
rect 70058 424170 78970 424226
rect 79026 424170 79094 424226
rect 79150 424170 79218 424226
rect 79274 424170 79342 424226
rect 79398 424170 96970 424226
rect 97026 424170 97094 424226
rect 97150 424170 97218 424226
rect 97274 424170 97342 424226
rect 97398 424170 100598 424226
rect 100654 424170 100722 424226
rect 100778 424170 131318 424226
rect 131374 424170 131442 424226
rect 131498 424170 162038 424226
rect 162094 424170 162162 424226
rect 162218 424170 192758 424226
rect 192814 424170 192882 424226
rect 192938 424170 223478 424226
rect 223534 424170 223602 424226
rect 223658 424170 254198 424226
rect 254254 424170 254322 424226
rect 254378 424170 284918 424226
rect 284974 424170 285042 424226
rect 285098 424170 315638 424226
rect 315694 424170 315762 424226
rect 315818 424170 346358 424226
rect 346414 424170 346482 424226
rect 346538 424170 377078 424226
rect 377134 424170 377202 424226
rect 377258 424170 407798 424226
rect 407854 424170 407922 424226
rect 407978 424170 438518 424226
rect 438574 424170 438642 424226
rect 438698 424170 469238 424226
rect 469294 424170 469362 424226
rect 469418 424170 499958 424226
rect 500014 424170 500082 424226
rect 500138 424170 530678 424226
rect 530734 424170 530802 424226
rect 530858 424170 564970 424226
rect 565026 424170 565094 424226
rect 565150 424170 565218 424226
rect 565274 424170 565342 424226
rect 565398 424170 582970 424226
rect 583026 424170 583094 424226
rect 583150 424170 583218 424226
rect 583274 424170 583342 424226
rect 583398 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect -1916 424102 597980 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 6970 424102
rect 7026 424046 7094 424102
rect 7150 424046 7218 424102
rect 7274 424046 7342 424102
rect 7398 424046 24970 424102
rect 25026 424046 25094 424102
rect 25150 424046 25218 424102
rect 25274 424046 25342 424102
rect 25398 424046 42970 424102
rect 43026 424046 43094 424102
rect 43150 424046 43218 424102
rect 43274 424046 43342 424102
rect 43398 424046 60970 424102
rect 61026 424046 61094 424102
rect 61150 424046 61218 424102
rect 61274 424046 61342 424102
rect 61398 424046 69878 424102
rect 69934 424046 70002 424102
rect 70058 424046 78970 424102
rect 79026 424046 79094 424102
rect 79150 424046 79218 424102
rect 79274 424046 79342 424102
rect 79398 424046 96970 424102
rect 97026 424046 97094 424102
rect 97150 424046 97218 424102
rect 97274 424046 97342 424102
rect 97398 424046 100598 424102
rect 100654 424046 100722 424102
rect 100778 424046 131318 424102
rect 131374 424046 131442 424102
rect 131498 424046 162038 424102
rect 162094 424046 162162 424102
rect 162218 424046 192758 424102
rect 192814 424046 192882 424102
rect 192938 424046 223478 424102
rect 223534 424046 223602 424102
rect 223658 424046 254198 424102
rect 254254 424046 254322 424102
rect 254378 424046 284918 424102
rect 284974 424046 285042 424102
rect 285098 424046 315638 424102
rect 315694 424046 315762 424102
rect 315818 424046 346358 424102
rect 346414 424046 346482 424102
rect 346538 424046 377078 424102
rect 377134 424046 377202 424102
rect 377258 424046 407798 424102
rect 407854 424046 407922 424102
rect 407978 424046 438518 424102
rect 438574 424046 438642 424102
rect 438698 424046 469238 424102
rect 469294 424046 469362 424102
rect 469418 424046 499958 424102
rect 500014 424046 500082 424102
rect 500138 424046 530678 424102
rect 530734 424046 530802 424102
rect 530858 424046 564970 424102
rect 565026 424046 565094 424102
rect 565150 424046 565218 424102
rect 565274 424046 565342 424102
rect 565398 424046 582970 424102
rect 583026 424046 583094 424102
rect 583150 424046 583218 424102
rect 583274 424046 583342 424102
rect 583398 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect -1916 423978 597980 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 6970 423978
rect 7026 423922 7094 423978
rect 7150 423922 7218 423978
rect 7274 423922 7342 423978
rect 7398 423922 24970 423978
rect 25026 423922 25094 423978
rect 25150 423922 25218 423978
rect 25274 423922 25342 423978
rect 25398 423922 42970 423978
rect 43026 423922 43094 423978
rect 43150 423922 43218 423978
rect 43274 423922 43342 423978
rect 43398 423922 60970 423978
rect 61026 423922 61094 423978
rect 61150 423922 61218 423978
rect 61274 423922 61342 423978
rect 61398 423922 69878 423978
rect 69934 423922 70002 423978
rect 70058 423922 78970 423978
rect 79026 423922 79094 423978
rect 79150 423922 79218 423978
rect 79274 423922 79342 423978
rect 79398 423922 96970 423978
rect 97026 423922 97094 423978
rect 97150 423922 97218 423978
rect 97274 423922 97342 423978
rect 97398 423922 100598 423978
rect 100654 423922 100722 423978
rect 100778 423922 131318 423978
rect 131374 423922 131442 423978
rect 131498 423922 162038 423978
rect 162094 423922 162162 423978
rect 162218 423922 192758 423978
rect 192814 423922 192882 423978
rect 192938 423922 223478 423978
rect 223534 423922 223602 423978
rect 223658 423922 254198 423978
rect 254254 423922 254322 423978
rect 254378 423922 284918 423978
rect 284974 423922 285042 423978
rect 285098 423922 315638 423978
rect 315694 423922 315762 423978
rect 315818 423922 346358 423978
rect 346414 423922 346482 423978
rect 346538 423922 377078 423978
rect 377134 423922 377202 423978
rect 377258 423922 407798 423978
rect 407854 423922 407922 423978
rect 407978 423922 438518 423978
rect 438574 423922 438642 423978
rect 438698 423922 469238 423978
rect 469294 423922 469362 423978
rect 469418 423922 499958 423978
rect 500014 423922 500082 423978
rect 500138 423922 530678 423978
rect 530734 423922 530802 423978
rect 530858 423922 564970 423978
rect 565026 423922 565094 423978
rect 565150 423922 565218 423978
rect 565274 423922 565342 423978
rect 565398 423922 582970 423978
rect 583026 423922 583094 423978
rect 583150 423922 583218 423978
rect 583274 423922 583342 423978
rect 583398 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect -1916 423826 597980 423922
rect -1916 418350 597980 418446
rect -1916 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 3250 418350
rect 3306 418294 3374 418350
rect 3430 418294 3498 418350
rect 3554 418294 3622 418350
rect 3678 418294 21250 418350
rect 21306 418294 21374 418350
rect 21430 418294 21498 418350
rect 21554 418294 21622 418350
rect 21678 418294 39250 418350
rect 39306 418294 39374 418350
rect 39430 418294 39498 418350
rect 39554 418294 39622 418350
rect 39678 418294 54518 418350
rect 54574 418294 54642 418350
rect 54698 418294 57250 418350
rect 57306 418294 57374 418350
rect 57430 418294 57498 418350
rect 57554 418294 57622 418350
rect 57678 418294 75250 418350
rect 75306 418294 75374 418350
rect 75430 418294 75498 418350
rect 75554 418294 75622 418350
rect 75678 418294 85238 418350
rect 85294 418294 85362 418350
rect 85418 418294 93250 418350
rect 93306 418294 93374 418350
rect 93430 418294 93498 418350
rect 93554 418294 93622 418350
rect 93678 418294 111250 418350
rect 111306 418294 111374 418350
rect 111430 418294 111498 418350
rect 111554 418294 111622 418350
rect 111678 418294 115958 418350
rect 116014 418294 116082 418350
rect 116138 418294 146678 418350
rect 146734 418294 146802 418350
rect 146858 418294 177398 418350
rect 177454 418294 177522 418350
rect 177578 418294 208118 418350
rect 208174 418294 208242 418350
rect 208298 418294 238838 418350
rect 238894 418294 238962 418350
rect 239018 418294 269558 418350
rect 269614 418294 269682 418350
rect 269738 418294 300278 418350
rect 300334 418294 300402 418350
rect 300458 418294 330998 418350
rect 331054 418294 331122 418350
rect 331178 418294 361718 418350
rect 361774 418294 361842 418350
rect 361898 418294 392438 418350
rect 392494 418294 392562 418350
rect 392618 418294 423158 418350
rect 423214 418294 423282 418350
rect 423338 418294 453878 418350
rect 453934 418294 454002 418350
rect 454058 418294 484598 418350
rect 484654 418294 484722 418350
rect 484778 418294 515318 418350
rect 515374 418294 515442 418350
rect 515498 418294 546038 418350
rect 546094 418294 546162 418350
rect 546218 418294 561250 418350
rect 561306 418294 561374 418350
rect 561430 418294 561498 418350
rect 561554 418294 561622 418350
rect 561678 418294 579250 418350
rect 579306 418294 579374 418350
rect 579430 418294 579498 418350
rect 579554 418294 579622 418350
rect 579678 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597980 418350
rect -1916 418226 597980 418294
rect -1916 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 3250 418226
rect 3306 418170 3374 418226
rect 3430 418170 3498 418226
rect 3554 418170 3622 418226
rect 3678 418170 21250 418226
rect 21306 418170 21374 418226
rect 21430 418170 21498 418226
rect 21554 418170 21622 418226
rect 21678 418170 39250 418226
rect 39306 418170 39374 418226
rect 39430 418170 39498 418226
rect 39554 418170 39622 418226
rect 39678 418170 54518 418226
rect 54574 418170 54642 418226
rect 54698 418170 57250 418226
rect 57306 418170 57374 418226
rect 57430 418170 57498 418226
rect 57554 418170 57622 418226
rect 57678 418170 75250 418226
rect 75306 418170 75374 418226
rect 75430 418170 75498 418226
rect 75554 418170 75622 418226
rect 75678 418170 85238 418226
rect 85294 418170 85362 418226
rect 85418 418170 93250 418226
rect 93306 418170 93374 418226
rect 93430 418170 93498 418226
rect 93554 418170 93622 418226
rect 93678 418170 111250 418226
rect 111306 418170 111374 418226
rect 111430 418170 111498 418226
rect 111554 418170 111622 418226
rect 111678 418170 115958 418226
rect 116014 418170 116082 418226
rect 116138 418170 146678 418226
rect 146734 418170 146802 418226
rect 146858 418170 177398 418226
rect 177454 418170 177522 418226
rect 177578 418170 208118 418226
rect 208174 418170 208242 418226
rect 208298 418170 238838 418226
rect 238894 418170 238962 418226
rect 239018 418170 269558 418226
rect 269614 418170 269682 418226
rect 269738 418170 300278 418226
rect 300334 418170 300402 418226
rect 300458 418170 330998 418226
rect 331054 418170 331122 418226
rect 331178 418170 361718 418226
rect 361774 418170 361842 418226
rect 361898 418170 392438 418226
rect 392494 418170 392562 418226
rect 392618 418170 423158 418226
rect 423214 418170 423282 418226
rect 423338 418170 453878 418226
rect 453934 418170 454002 418226
rect 454058 418170 484598 418226
rect 484654 418170 484722 418226
rect 484778 418170 515318 418226
rect 515374 418170 515442 418226
rect 515498 418170 546038 418226
rect 546094 418170 546162 418226
rect 546218 418170 561250 418226
rect 561306 418170 561374 418226
rect 561430 418170 561498 418226
rect 561554 418170 561622 418226
rect 561678 418170 579250 418226
rect 579306 418170 579374 418226
rect 579430 418170 579498 418226
rect 579554 418170 579622 418226
rect 579678 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597980 418226
rect -1916 418102 597980 418170
rect -1916 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 3250 418102
rect 3306 418046 3374 418102
rect 3430 418046 3498 418102
rect 3554 418046 3622 418102
rect 3678 418046 21250 418102
rect 21306 418046 21374 418102
rect 21430 418046 21498 418102
rect 21554 418046 21622 418102
rect 21678 418046 39250 418102
rect 39306 418046 39374 418102
rect 39430 418046 39498 418102
rect 39554 418046 39622 418102
rect 39678 418046 54518 418102
rect 54574 418046 54642 418102
rect 54698 418046 57250 418102
rect 57306 418046 57374 418102
rect 57430 418046 57498 418102
rect 57554 418046 57622 418102
rect 57678 418046 75250 418102
rect 75306 418046 75374 418102
rect 75430 418046 75498 418102
rect 75554 418046 75622 418102
rect 75678 418046 85238 418102
rect 85294 418046 85362 418102
rect 85418 418046 93250 418102
rect 93306 418046 93374 418102
rect 93430 418046 93498 418102
rect 93554 418046 93622 418102
rect 93678 418046 111250 418102
rect 111306 418046 111374 418102
rect 111430 418046 111498 418102
rect 111554 418046 111622 418102
rect 111678 418046 115958 418102
rect 116014 418046 116082 418102
rect 116138 418046 146678 418102
rect 146734 418046 146802 418102
rect 146858 418046 177398 418102
rect 177454 418046 177522 418102
rect 177578 418046 208118 418102
rect 208174 418046 208242 418102
rect 208298 418046 238838 418102
rect 238894 418046 238962 418102
rect 239018 418046 269558 418102
rect 269614 418046 269682 418102
rect 269738 418046 300278 418102
rect 300334 418046 300402 418102
rect 300458 418046 330998 418102
rect 331054 418046 331122 418102
rect 331178 418046 361718 418102
rect 361774 418046 361842 418102
rect 361898 418046 392438 418102
rect 392494 418046 392562 418102
rect 392618 418046 423158 418102
rect 423214 418046 423282 418102
rect 423338 418046 453878 418102
rect 453934 418046 454002 418102
rect 454058 418046 484598 418102
rect 484654 418046 484722 418102
rect 484778 418046 515318 418102
rect 515374 418046 515442 418102
rect 515498 418046 546038 418102
rect 546094 418046 546162 418102
rect 546218 418046 561250 418102
rect 561306 418046 561374 418102
rect 561430 418046 561498 418102
rect 561554 418046 561622 418102
rect 561678 418046 579250 418102
rect 579306 418046 579374 418102
rect 579430 418046 579498 418102
rect 579554 418046 579622 418102
rect 579678 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597980 418102
rect -1916 417978 597980 418046
rect -1916 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 3250 417978
rect 3306 417922 3374 417978
rect 3430 417922 3498 417978
rect 3554 417922 3622 417978
rect 3678 417922 21250 417978
rect 21306 417922 21374 417978
rect 21430 417922 21498 417978
rect 21554 417922 21622 417978
rect 21678 417922 39250 417978
rect 39306 417922 39374 417978
rect 39430 417922 39498 417978
rect 39554 417922 39622 417978
rect 39678 417922 54518 417978
rect 54574 417922 54642 417978
rect 54698 417922 57250 417978
rect 57306 417922 57374 417978
rect 57430 417922 57498 417978
rect 57554 417922 57622 417978
rect 57678 417922 75250 417978
rect 75306 417922 75374 417978
rect 75430 417922 75498 417978
rect 75554 417922 75622 417978
rect 75678 417922 85238 417978
rect 85294 417922 85362 417978
rect 85418 417922 93250 417978
rect 93306 417922 93374 417978
rect 93430 417922 93498 417978
rect 93554 417922 93622 417978
rect 93678 417922 111250 417978
rect 111306 417922 111374 417978
rect 111430 417922 111498 417978
rect 111554 417922 111622 417978
rect 111678 417922 115958 417978
rect 116014 417922 116082 417978
rect 116138 417922 146678 417978
rect 146734 417922 146802 417978
rect 146858 417922 177398 417978
rect 177454 417922 177522 417978
rect 177578 417922 208118 417978
rect 208174 417922 208242 417978
rect 208298 417922 238838 417978
rect 238894 417922 238962 417978
rect 239018 417922 269558 417978
rect 269614 417922 269682 417978
rect 269738 417922 300278 417978
rect 300334 417922 300402 417978
rect 300458 417922 330998 417978
rect 331054 417922 331122 417978
rect 331178 417922 361718 417978
rect 361774 417922 361842 417978
rect 361898 417922 392438 417978
rect 392494 417922 392562 417978
rect 392618 417922 423158 417978
rect 423214 417922 423282 417978
rect 423338 417922 453878 417978
rect 453934 417922 454002 417978
rect 454058 417922 484598 417978
rect 484654 417922 484722 417978
rect 484778 417922 515318 417978
rect 515374 417922 515442 417978
rect 515498 417922 546038 417978
rect 546094 417922 546162 417978
rect 546218 417922 561250 417978
rect 561306 417922 561374 417978
rect 561430 417922 561498 417978
rect 561554 417922 561622 417978
rect 561678 417922 579250 417978
rect 579306 417922 579374 417978
rect 579430 417922 579498 417978
rect 579554 417922 579622 417978
rect 579678 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597980 417978
rect -1916 417826 597980 417922
rect -1916 406350 597980 406446
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 6970 406350
rect 7026 406294 7094 406350
rect 7150 406294 7218 406350
rect 7274 406294 7342 406350
rect 7398 406294 24970 406350
rect 25026 406294 25094 406350
rect 25150 406294 25218 406350
rect 25274 406294 25342 406350
rect 25398 406294 42970 406350
rect 43026 406294 43094 406350
rect 43150 406294 43218 406350
rect 43274 406294 43342 406350
rect 43398 406294 60970 406350
rect 61026 406294 61094 406350
rect 61150 406294 61218 406350
rect 61274 406294 61342 406350
rect 61398 406294 69878 406350
rect 69934 406294 70002 406350
rect 70058 406294 78970 406350
rect 79026 406294 79094 406350
rect 79150 406294 79218 406350
rect 79274 406294 79342 406350
rect 79398 406294 96970 406350
rect 97026 406294 97094 406350
rect 97150 406294 97218 406350
rect 97274 406294 97342 406350
rect 97398 406294 100598 406350
rect 100654 406294 100722 406350
rect 100778 406294 131318 406350
rect 131374 406294 131442 406350
rect 131498 406294 162038 406350
rect 162094 406294 162162 406350
rect 162218 406294 192758 406350
rect 192814 406294 192882 406350
rect 192938 406294 223478 406350
rect 223534 406294 223602 406350
rect 223658 406294 254198 406350
rect 254254 406294 254322 406350
rect 254378 406294 284918 406350
rect 284974 406294 285042 406350
rect 285098 406294 315638 406350
rect 315694 406294 315762 406350
rect 315818 406294 346358 406350
rect 346414 406294 346482 406350
rect 346538 406294 377078 406350
rect 377134 406294 377202 406350
rect 377258 406294 407798 406350
rect 407854 406294 407922 406350
rect 407978 406294 438518 406350
rect 438574 406294 438642 406350
rect 438698 406294 469238 406350
rect 469294 406294 469362 406350
rect 469418 406294 499958 406350
rect 500014 406294 500082 406350
rect 500138 406294 530678 406350
rect 530734 406294 530802 406350
rect 530858 406294 564970 406350
rect 565026 406294 565094 406350
rect 565150 406294 565218 406350
rect 565274 406294 565342 406350
rect 565398 406294 582970 406350
rect 583026 406294 583094 406350
rect 583150 406294 583218 406350
rect 583274 406294 583342 406350
rect 583398 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect -1916 406226 597980 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 6970 406226
rect 7026 406170 7094 406226
rect 7150 406170 7218 406226
rect 7274 406170 7342 406226
rect 7398 406170 24970 406226
rect 25026 406170 25094 406226
rect 25150 406170 25218 406226
rect 25274 406170 25342 406226
rect 25398 406170 42970 406226
rect 43026 406170 43094 406226
rect 43150 406170 43218 406226
rect 43274 406170 43342 406226
rect 43398 406170 60970 406226
rect 61026 406170 61094 406226
rect 61150 406170 61218 406226
rect 61274 406170 61342 406226
rect 61398 406170 69878 406226
rect 69934 406170 70002 406226
rect 70058 406170 78970 406226
rect 79026 406170 79094 406226
rect 79150 406170 79218 406226
rect 79274 406170 79342 406226
rect 79398 406170 96970 406226
rect 97026 406170 97094 406226
rect 97150 406170 97218 406226
rect 97274 406170 97342 406226
rect 97398 406170 100598 406226
rect 100654 406170 100722 406226
rect 100778 406170 131318 406226
rect 131374 406170 131442 406226
rect 131498 406170 162038 406226
rect 162094 406170 162162 406226
rect 162218 406170 192758 406226
rect 192814 406170 192882 406226
rect 192938 406170 223478 406226
rect 223534 406170 223602 406226
rect 223658 406170 254198 406226
rect 254254 406170 254322 406226
rect 254378 406170 284918 406226
rect 284974 406170 285042 406226
rect 285098 406170 315638 406226
rect 315694 406170 315762 406226
rect 315818 406170 346358 406226
rect 346414 406170 346482 406226
rect 346538 406170 377078 406226
rect 377134 406170 377202 406226
rect 377258 406170 407798 406226
rect 407854 406170 407922 406226
rect 407978 406170 438518 406226
rect 438574 406170 438642 406226
rect 438698 406170 469238 406226
rect 469294 406170 469362 406226
rect 469418 406170 499958 406226
rect 500014 406170 500082 406226
rect 500138 406170 530678 406226
rect 530734 406170 530802 406226
rect 530858 406170 564970 406226
rect 565026 406170 565094 406226
rect 565150 406170 565218 406226
rect 565274 406170 565342 406226
rect 565398 406170 582970 406226
rect 583026 406170 583094 406226
rect 583150 406170 583218 406226
rect 583274 406170 583342 406226
rect 583398 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect -1916 406102 597980 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 6970 406102
rect 7026 406046 7094 406102
rect 7150 406046 7218 406102
rect 7274 406046 7342 406102
rect 7398 406046 24970 406102
rect 25026 406046 25094 406102
rect 25150 406046 25218 406102
rect 25274 406046 25342 406102
rect 25398 406046 42970 406102
rect 43026 406046 43094 406102
rect 43150 406046 43218 406102
rect 43274 406046 43342 406102
rect 43398 406046 60970 406102
rect 61026 406046 61094 406102
rect 61150 406046 61218 406102
rect 61274 406046 61342 406102
rect 61398 406046 69878 406102
rect 69934 406046 70002 406102
rect 70058 406046 78970 406102
rect 79026 406046 79094 406102
rect 79150 406046 79218 406102
rect 79274 406046 79342 406102
rect 79398 406046 96970 406102
rect 97026 406046 97094 406102
rect 97150 406046 97218 406102
rect 97274 406046 97342 406102
rect 97398 406046 100598 406102
rect 100654 406046 100722 406102
rect 100778 406046 131318 406102
rect 131374 406046 131442 406102
rect 131498 406046 162038 406102
rect 162094 406046 162162 406102
rect 162218 406046 192758 406102
rect 192814 406046 192882 406102
rect 192938 406046 223478 406102
rect 223534 406046 223602 406102
rect 223658 406046 254198 406102
rect 254254 406046 254322 406102
rect 254378 406046 284918 406102
rect 284974 406046 285042 406102
rect 285098 406046 315638 406102
rect 315694 406046 315762 406102
rect 315818 406046 346358 406102
rect 346414 406046 346482 406102
rect 346538 406046 377078 406102
rect 377134 406046 377202 406102
rect 377258 406046 407798 406102
rect 407854 406046 407922 406102
rect 407978 406046 438518 406102
rect 438574 406046 438642 406102
rect 438698 406046 469238 406102
rect 469294 406046 469362 406102
rect 469418 406046 499958 406102
rect 500014 406046 500082 406102
rect 500138 406046 530678 406102
rect 530734 406046 530802 406102
rect 530858 406046 564970 406102
rect 565026 406046 565094 406102
rect 565150 406046 565218 406102
rect 565274 406046 565342 406102
rect 565398 406046 582970 406102
rect 583026 406046 583094 406102
rect 583150 406046 583218 406102
rect 583274 406046 583342 406102
rect 583398 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect -1916 405978 597980 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 6970 405978
rect 7026 405922 7094 405978
rect 7150 405922 7218 405978
rect 7274 405922 7342 405978
rect 7398 405922 24970 405978
rect 25026 405922 25094 405978
rect 25150 405922 25218 405978
rect 25274 405922 25342 405978
rect 25398 405922 42970 405978
rect 43026 405922 43094 405978
rect 43150 405922 43218 405978
rect 43274 405922 43342 405978
rect 43398 405922 60970 405978
rect 61026 405922 61094 405978
rect 61150 405922 61218 405978
rect 61274 405922 61342 405978
rect 61398 405922 69878 405978
rect 69934 405922 70002 405978
rect 70058 405922 78970 405978
rect 79026 405922 79094 405978
rect 79150 405922 79218 405978
rect 79274 405922 79342 405978
rect 79398 405922 96970 405978
rect 97026 405922 97094 405978
rect 97150 405922 97218 405978
rect 97274 405922 97342 405978
rect 97398 405922 100598 405978
rect 100654 405922 100722 405978
rect 100778 405922 131318 405978
rect 131374 405922 131442 405978
rect 131498 405922 162038 405978
rect 162094 405922 162162 405978
rect 162218 405922 192758 405978
rect 192814 405922 192882 405978
rect 192938 405922 223478 405978
rect 223534 405922 223602 405978
rect 223658 405922 254198 405978
rect 254254 405922 254322 405978
rect 254378 405922 284918 405978
rect 284974 405922 285042 405978
rect 285098 405922 315638 405978
rect 315694 405922 315762 405978
rect 315818 405922 346358 405978
rect 346414 405922 346482 405978
rect 346538 405922 377078 405978
rect 377134 405922 377202 405978
rect 377258 405922 407798 405978
rect 407854 405922 407922 405978
rect 407978 405922 438518 405978
rect 438574 405922 438642 405978
rect 438698 405922 469238 405978
rect 469294 405922 469362 405978
rect 469418 405922 499958 405978
rect 500014 405922 500082 405978
rect 500138 405922 530678 405978
rect 530734 405922 530802 405978
rect 530858 405922 564970 405978
rect 565026 405922 565094 405978
rect 565150 405922 565218 405978
rect 565274 405922 565342 405978
rect 565398 405922 582970 405978
rect 583026 405922 583094 405978
rect 583150 405922 583218 405978
rect 583274 405922 583342 405978
rect 583398 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect -1916 405826 597980 405922
rect -1916 400350 597980 400446
rect -1916 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 3250 400350
rect 3306 400294 3374 400350
rect 3430 400294 3498 400350
rect 3554 400294 3622 400350
rect 3678 400294 21250 400350
rect 21306 400294 21374 400350
rect 21430 400294 21498 400350
rect 21554 400294 21622 400350
rect 21678 400294 39250 400350
rect 39306 400294 39374 400350
rect 39430 400294 39498 400350
rect 39554 400294 39622 400350
rect 39678 400294 54518 400350
rect 54574 400294 54642 400350
rect 54698 400294 57250 400350
rect 57306 400294 57374 400350
rect 57430 400294 57498 400350
rect 57554 400294 57622 400350
rect 57678 400294 75250 400350
rect 75306 400294 75374 400350
rect 75430 400294 75498 400350
rect 75554 400294 75622 400350
rect 75678 400294 85238 400350
rect 85294 400294 85362 400350
rect 85418 400294 93250 400350
rect 93306 400294 93374 400350
rect 93430 400294 93498 400350
rect 93554 400294 93622 400350
rect 93678 400294 111250 400350
rect 111306 400294 111374 400350
rect 111430 400294 111498 400350
rect 111554 400294 111622 400350
rect 111678 400294 115958 400350
rect 116014 400294 116082 400350
rect 116138 400294 146678 400350
rect 146734 400294 146802 400350
rect 146858 400294 177398 400350
rect 177454 400294 177522 400350
rect 177578 400294 208118 400350
rect 208174 400294 208242 400350
rect 208298 400294 238838 400350
rect 238894 400294 238962 400350
rect 239018 400294 269558 400350
rect 269614 400294 269682 400350
rect 269738 400294 300278 400350
rect 300334 400294 300402 400350
rect 300458 400294 330998 400350
rect 331054 400294 331122 400350
rect 331178 400294 361718 400350
rect 361774 400294 361842 400350
rect 361898 400294 392438 400350
rect 392494 400294 392562 400350
rect 392618 400294 423158 400350
rect 423214 400294 423282 400350
rect 423338 400294 453878 400350
rect 453934 400294 454002 400350
rect 454058 400294 484598 400350
rect 484654 400294 484722 400350
rect 484778 400294 515318 400350
rect 515374 400294 515442 400350
rect 515498 400294 546038 400350
rect 546094 400294 546162 400350
rect 546218 400294 561250 400350
rect 561306 400294 561374 400350
rect 561430 400294 561498 400350
rect 561554 400294 561622 400350
rect 561678 400294 579250 400350
rect 579306 400294 579374 400350
rect 579430 400294 579498 400350
rect 579554 400294 579622 400350
rect 579678 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597980 400350
rect -1916 400226 597980 400294
rect -1916 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 3250 400226
rect 3306 400170 3374 400226
rect 3430 400170 3498 400226
rect 3554 400170 3622 400226
rect 3678 400170 21250 400226
rect 21306 400170 21374 400226
rect 21430 400170 21498 400226
rect 21554 400170 21622 400226
rect 21678 400170 39250 400226
rect 39306 400170 39374 400226
rect 39430 400170 39498 400226
rect 39554 400170 39622 400226
rect 39678 400170 54518 400226
rect 54574 400170 54642 400226
rect 54698 400170 57250 400226
rect 57306 400170 57374 400226
rect 57430 400170 57498 400226
rect 57554 400170 57622 400226
rect 57678 400170 75250 400226
rect 75306 400170 75374 400226
rect 75430 400170 75498 400226
rect 75554 400170 75622 400226
rect 75678 400170 85238 400226
rect 85294 400170 85362 400226
rect 85418 400170 93250 400226
rect 93306 400170 93374 400226
rect 93430 400170 93498 400226
rect 93554 400170 93622 400226
rect 93678 400170 111250 400226
rect 111306 400170 111374 400226
rect 111430 400170 111498 400226
rect 111554 400170 111622 400226
rect 111678 400170 115958 400226
rect 116014 400170 116082 400226
rect 116138 400170 146678 400226
rect 146734 400170 146802 400226
rect 146858 400170 177398 400226
rect 177454 400170 177522 400226
rect 177578 400170 208118 400226
rect 208174 400170 208242 400226
rect 208298 400170 238838 400226
rect 238894 400170 238962 400226
rect 239018 400170 269558 400226
rect 269614 400170 269682 400226
rect 269738 400170 300278 400226
rect 300334 400170 300402 400226
rect 300458 400170 330998 400226
rect 331054 400170 331122 400226
rect 331178 400170 361718 400226
rect 361774 400170 361842 400226
rect 361898 400170 392438 400226
rect 392494 400170 392562 400226
rect 392618 400170 423158 400226
rect 423214 400170 423282 400226
rect 423338 400170 453878 400226
rect 453934 400170 454002 400226
rect 454058 400170 484598 400226
rect 484654 400170 484722 400226
rect 484778 400170 515318 400226
rect 515374 400170 515442 400226
rect 515498 400170 546038 400226
rect 546094 400170 546162 400226
rect 546218 400170 561250 400226
rect 561306 400170 561374 400226
rect 561430 400170 561498 400226
rect 561554 400170 561622 400226
rect 561678 400170 579250 400226
rect 579306 400170 579374 400226
rect 579430 400170 579498 400226
rect 579554 400170 579622 400226
rect 579678 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597980 400226
rect -1916 400102 597980 400170
rect -1916 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 3250 400102
rect 3306 400046 3374 400102
rect 3430 400046 3498 400102
rect 3554 400046 3622 400102
rect 3678 400046 21250 400102
rect 21306 400046 21374 400102
rect 21430 400046 21498 400102
rect 21554 400046 21622 400102
rect 21678 400046 39250 400102
rect 39306 400046 39374 400102
rect 39430 400046 39498 400102
rect 39554 400046 39622 400102
rect 39678 400046 54518 400102
rect 54574 400046 54642 400102
rect 54698 400046 57250 400102
rect 57306 400046 57374 400102
rect 57430 400046 57498 400102
rect 57554 400046 57622 400102
rect 57678 400046 75250 400102
rect 75306 400046 75374 400102
rect 75430 400046 75498 400102
rect 75554 400046 75622 400102
rect 75678 400046 85238 400102
rect 85294 400046 85362 400102
rect 85418 400046 93250 400102
rect 93306 400046 93374 400102
rect 93430 400046 93498 400102
rect 93554 400046 93622 400102
rect 93678 400046 111250 400102
rect 111306 400046 111374 400102
rect 111430 400046 111498 400102
rect 111554 400046 111622 400102
rect 111678 400046 115958 400102
rect 116014 400046 116082 400102
rect 116138 400046 146678 400102
rect 146734 400046 146802 400102
rect 146858 400046 177398 400102
rect 177454 400046 177522 400102
rect 177578 400046 208118 400102
rect 208174 400046 208242 400102
rect 208298 400046 238838 400102
rect 238894 400046 238962 400102
rect 239018 400046 269558 400102
rect 269614 400046 269682 400102
rect 269738 400046 300278 400102
rect 300334 400046 300402 400102
rect 300458 400046 330998 400102
rect 331054 400046 331122 400102
rect 331178 400046 361718 400102
rect 361774 400046 361842 400102
rect 361898 400046 392438 400102
rect 392494 400046 392562 400102
rect 392618 400046 423158 400102
rect 423214 400046 423282 400102
rect 423338 400046 453878 400102
rect 453934 400046 454002 400102
rect 454058 400046 484598 400102
rect 484654 400046 484722 400102
rect 484778 400046 515318 400102
rect 515374 400046 515442 400102
rect 515498 400046 546038 400102
rect 546094 400046 546162 400102
rect 546218 400046 561250 400102
rect 561306 400046 561374 400102
rect 561430 400046 561498 400102
rect 561554 400046 561622 400102
rect 561678 400046 579250 400102
rect 579306 400046 579374 400102
rect 579430 400046 579498 400102
rect 579554 400046 579622 400102
rect 579678 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597980 400102
rect -1916 399978 597980 400046
rect -1916 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 3250 399978
rect 3306 399922 3374 399978
rect 3430 399922 3498 399978
rect 3554 399922 3622 399978
rect 3678 399922 21250 399978
rect 21306 399922 21374 399978
rect 21430 399922 21498 399978
rect 21554 399922 21622 399978
rect 21678 399922 39250 399978
rect 39306 399922 39374 399978
rect 39430 399922 39498 399978
rect 39554 399922 39622 399978
rect 39678 399922 54518 399978
rect 54574 399922 54642 399978
rect 54698 399922 57250 399978
rect 57306 399922 57374 399978
rect 57430 399922 57498 399978
rect 57554 399922 57622 399978
rect 57678 399922 75250 399978
rect 75306 399922 75374 399978
rect 75430 399922 75498 399978
rect 75554 399922 75622 399978
rect 75678 399922 85238 399978
rect 85294 399922 85362 399978
rect 85418 399922 93250 399978
rect 93306 399922 93374 399978
rect 93430 399922 93498 399978
rect 93554 399922 93622 399978
rect 93678 399922 111250 399978
rect 111306 399922 111374 399978
rect 111430 399922 111498 399978
rect 111554 399922 111622 399978
rect 111678 399922 115958 399978
rect 116014 399922 116082 399978
rect 116138 399922 146678 399978
rect 146734 399922 146802 399978
rect 146858 399922 177398 399978
rect 177454 399922 177522 399978
rect 177578 399922 208118 399978
rect 208174 399922 208242 399978
rect 208298 399922 238838 399978
rect 238894 399922 238962 399978
rect 239018 399922 269558 399978
rect 269614 399922 269682 399978
rect 269738 399922 300278 399978
rect 300334 399922 300402 399978
rect 300458 399922 330998 399978
rect 331054 399922 331122 399978
rect 331178 399922 361718 399978
rect 361774 399922 361842 399978
rect 361898 399922 392438 399978
rect 392494 399922 392562 399978
rect 392618 399922 423158 399978
rect 423214 399922 423282 399978
rect 423338 399922 453878 399978
rect 453934 399922 454002 399978
rect 454058 399922 484598 399978
rect 484654 399922 484722 399978
rect 484778 399922 515318 399978
rect 515374 399922 515442 399978
rect 515498 399922 546038 399978
rect 546094 399922 546162 399978
rect 546218 399922 561250 399978
rect 561306 399922 561374 399978
rect 561430 399922 561498 399978
rect 561554 399922 561622 399978
rect 561678 399922 579250 399978
rect 579306 399922 579374 399978
rect 579430 399922 579498 399978
rect 579554 399922 579622 399978
rect 579678 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597980 399978
rect -1916 399826 597980 399922
rect -1916 388350 597980 388446
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 6970 388350
rect 7026 388294 7094 388350
rect 7150 388294 7218 388350
rect 7274 388294 7342 388350
rect 7398 388294 24970 388350
rect 25026 388294 25094 388350
rect 25150 388294 25218 388350
rect 25274 388294 25342 388350
rect 25398 388294 42970 388350
rect 43026 388294 43094 388350
rect 43150 388294 43218 388350
rect 43274 388294 43342 388350
rect 43398 388294 60970 388350
rect 61026 388294 61094 388350
rect 61150 388294 61218 388350
rect 61274 388294 61342 388350
rect 61398 388294 69878 388350
rect 69934 388294 70002 388350
rect 70058 388294 78970 388350
rect 79026 388294 79094 388350
rect 79150 388294 79218 388350
rect 79274 388294 79342 388350
rect 79398 388294 96970 388350
rect 97026 388294 97094 388350
rect 97150 388294 97218 388350
rect 97274 388294 97342 388350
rect 97398 388294 100598 388350
rect 100654 388294 100722 388350
rect 100778 388294 131318 388350
rect 131374 388294 131442 388350
rect 131498 388294 162038 388350
rect 162094 388294 162162 388350
rect 162218 388294 192758 388350
rect 192814 388294 192882 388350
rect 192938 388294 223478 388350
rect 223534 388294 223602 388350
rect 223658 388294 254198 388350
rect 254254 388294 254322 388350
rect 254378 388294 284918 388350
rect 284974 388294 285042 388350
rect 285098 388294 315638 388350
rect 315694 388294 315762 388350
rect 315818 388294 346358 388350
rect 346414 388294 346482 388350
rect 346538 388294 377078 388350
rect 377134 388294 377202 388350
rect 377258 388294 407798 388350
rect 407854 388294 407922 388350
rect 407978 388294 438518 388350
rect 438574 388294 438642 388350
rect 438698 388294 469238 388350
rect 469294 388294 469362 388350
rect 469418 388294 499958 388350
rect 500014 388294 500082 388350
rect 500138 388294 530678 388350
rect 530734 388294 530802 388350
rect 530858 388294 564970 388350
rect 565026 388294 565094 388350
rect 565150 388294 565218 388350
rect 565274 388294 565342 388350
rect 565398 388294 582970 388350
rect 583026 388294 583094 388350
rect 583150 388294 583218 388350
rect 583274 388294 583342 388350
rect 583398 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect -1916 388226 597980 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 6970 388226
rect 7026 388170 7094 388226
rect 7150 388170 7218 388226
rect 7274 388170 7342 388226
rect 7398 388170 24970 388226
rect 25026 388170 25094 388226
rect 25150 388170 25218 388226
rect 25274 388170 25342 388226
rect 25398 388170 42970 388226
rect 43026 388170 43094 388226
rect 43150 388170 43218 388226
rect 43274 388170 43342 388226
rect 43398 388170 60970 388226
rect 61026 388170 61094 388226
rect 61150 388170 61218 388226
rect 61274 388170 61342 388226
rect 61398 388170 69878 388226
rect 69934 388170 70002 388226
rect 70058 388170 78970 388226
rect 79026 388170 79094 388226
rect 79150 388170 79218 388226
rect 79274 388170 79342 388226
rect 79398 388170 96970 388226
rect 97026 388170 97094 388226
rect 97150 388170 97218 388226
rect 97274 388170 97342 388226
rect 97398 388170 100598 388226
rect 100654 388170 100722 388226
rect 100778 388170 131318 388226
rect 131374 388170 131442 388226
rect 131498 388170 162038 388226
rect 162094 388170 162162 388226
rect 162218 388170 192758 388226
rect 192814 388170 192882 388226
rect 192938 388170 223478 388226
rect 223534 388170 223602 388226
rect 223658 388170 254198 388226
rect 254254 388170 254322 388226
rect 254378 388170 284918 388226
rect 284974 388170 285042 388226
rect 285098 388170 315638 388226
rect 315694 388170 315762 388226
rect 315818 388170 346358 388226
rect 346414 388170 346482 388226
rect 346538 388170 377078 388226
rect 377134 388170 377202 388226
rect 377258 388170 407798 388226
rect 407854 388170 407922 388226
rect 407978 388170 438518 388226
rect 438574 388170 438642 388226
rect 438698 388170 469238 388226
rect 469294 388170 469362 388226
rect 469418 388170 499958 388226
rect 500014 388170 500082 388226
rect 500138 388170 530678 388226
rect 530734 388170 530802 388226
rect 530858 388170 564970 388226
rect 565026 388170 565094 388226
rect 565150 388170 565218 388226
rect 565274 388170 565342 388226
rect 565398 388170 582970 388226
rect 583026 388170 583094 388226
rect 583150 388170 583218 388226
rect 583274 388170 583342 388226
rect 583398 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect -1916 388102 597980 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 6970 388102
rect 7026 388046 7094 388102
rect 7150 388046 7218 388102
rect 7274 388046 7342 388102
rect 7398 388046 24970 388102
rect 25026 388046 25094 388102
rect 25150 388046 25218 388102
rect 25274 388046 25342 388102
rect 25398 388046 42970 388102
rect 43026 388046 43094 388102
rect 43150 388046 43218 388102
rect 43274 388046 43342 388102
rect 43398 388046 60970 388102
rect 61026 388046 61094 388102
rect 61150 388046 61218 388102
rect 61274 388046 61342 388102
rect 61398 388046 69878 388102
rect 69934 388046 70002 388102
rect 70058 388046 78970 388102
rect 79026 388046 79094 388102
rect 79150 388046 79218 388102
rect 79274 388046 79342 388102
rect 79398 388046 96970 388102
rect 97026 388046 97094 388102
rect 97150 388046 97218 388102
rect 97274 388046 97342 388102
rect 97398 388046 100598 388102
rect 100654 388046 100722 388102
rect 100778 388046 131318 388102
rect 131374 388046 131442 388102
rect 131498 388046 162038 388102
rect 162094 388046 162162 388102
rect 162218 388046 192758 388102
rect 192814 388046 192882 388102
rect 192938 388046 223478 388102
rect 223534 388046 223602 388102
rect 223658 388046 254198 388102
rect 254254 388046 254322 388102
rect 254378 388046 284918 388102
rect 284974 388046 285042 388102
rect 285098 388046 315638 388102
rect 315694 388046 315762 388102
rect 315818 388046 346358 388102
rect 346414 388046 346482 388102
rect 346538 388046 377078 388102
rect 377134 388046 377202 388102
rect 377258 388046 407798 388102
rect 407854 388046 407922 388102
rect 407978 388046 438518 388102
rect 438574 388046 438642 388102
rect 438698 388046 469238 388102
rect 469294 388046 469362 388102
rect 469418 388046 499958 388102
rect 500014 388046 500082 388102
rect 500138 388046 530678 388102
rect 530734 388046 530802 388102
rect 530858 388046 564970 388102
rect 565026 388046 565094 388102
rect 565150 388046 565218 388102
rect 565274 388046 565342 388102
rect 565398 388046 582970 388102
rect 583026 388046 583094 388102
rect 583150 388046 583218 388102
rect 583274 388046 583342 388102
rect 583398 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect -1916 387978 597980 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 6970 387978
rect 7026 387922 7094 387978
rect 7150 387922 7218 387978
rect 7274 387922 7342 387978
rect 7398 387922 24970 387978
rect 25026 387922 25094 387978
rect 25150 387922 25218 387978
rect 25274 387922 25342 387978
rect 25398 387922 42970 387978
rect 43026 387922 43094 387978
rect 43150 387922 43218 387978
rect 43274 387922 43342 387978
rect 43398 387922 60970 387978
rect 61026 387922 61094 387978
rect 61150 387922 61218 387978
rect 61274 387922 61342 387978
rect 61398 387922 69878 387978
rect 69934 387922 70002 387978
rect 70058 387922 78970 387978
rect 79026 387922 79094 387978
rect 79150 387922 79218 387978
rect 79274 387922 79342 387978
rect 79398 387922 96970 387978
rect 97026 387922 97094 387978
rect 97150 387922 97218 387978
rect 97274 387922 97342 387978
rect 97398 387922 100598 387978
rect 100654 387922 100722 387978
rect 100778 387922 131318 387978
rect 131374 387922 131442 387978
rect 131498 387922 162038 387978
rect 162094 387922 162162 387978
rect 162218 387922 192758 387978
rect 192814 387922 192882 387978
rect 192938 387922 223478 387978
rect 223534 387922 223602 387978
rect 223658 387922 254198 387978
rect 254254 387922 254322 387978
rect 254378 387922 284918 387978
rect 284974 387922 285042 387978
rect 285098 387922 315638 387978
rect 315694 387922 315762 387978
rect 315818 387922 346358 387978
rect 346414 387922 346482 387978
rect 346538 387922 377078 387978
rect 377134 387922 377202 387978
rect 377258 387922 407798 387978
rect 407854 387922 407922 387978
rect 407978 387922 438518 387978
rect 438574 387922 438642 387978
rect 438698 387922 469238 387978
rect 469294 387922 469362 387978
rect 469418 387922 499958 387978
rect 500014 387922 500082 387978
rect 500138 387922 530678 387978
rect 530734 387922 530802 387978
rect 530858 387922 564970 387978
rect 565026 387922 565094 387978
rect 565150 387922 565218 387978
rect 565274 387922 565342 387978
rect 565398 387922 582970 387978
rect 583026 387922 583094 387978
rect 583150 387922 583218 387978
rect 583274 387922 583342 387978
rect 583398 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect -1916 387826 597980 387922
rect -1916 382350 597980 382446
rect -1916 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 3250 382350
rect 3306 382294 3374 382350
rect 3430 382294 3498 382350
rect 3554 382294 3622 382350
rect 3678 382294 21250 382350
rect 21306 382294 21374 382350
rect 21430 382294 21498 382350
rect 21554 382294 21622 382350
rect 21678 382294 39250 382350
rect 39306 382294 39374 382350
rect 39430 382294 39498 382350
rect 39554 382294 39622 382350
rect 39678 382294 54518 382350
rect 54574 382294 54642 382350
rect 54698 382294 57250 382350
rect 57306 382294 57374 382350
rect 57430 382294 57498 382350
rect 57554 382294 57622 382350
rect 57678 382294 75250 382350
rect 75306 382294 75374 382350
rect 75430 382294 75498 382350
rect 75554 382294 75622 382350
rect 75678 382294 85238 382350
rect 85294 382294 85362 382350
rect 85418 382294 93250 382350
rect 93306 382294 93374 382350
rect 93430 382294 93498 382350
rect 93554 382294 93622 382350
rect 93678 382294 111250 382350
rect 111306 382294 111374 382350
rect 111430 382294 111498 382350
rect 111554 382294 111622 382350
rect 111678 382294 115958 382350
rect 116014 382294 116082 382350
rect 116138 382294 146678 382350
rect 146734 382294 146802 382350
rect 146858 382294 177398 382350
rect 177454 382294 177522 382350
rect 177578 382294 208118 382350
rect 208174 382294 208242 382350
rect 208298 382294 238838 382350
rect 238894 382294 238962 382350
rect 239018 382294 269558 382350
rect 269614 382294 269682 382350
rect 269738 382294 300278 382350
rect 300334 382294 300402 382350
rect 300458 382294 330998 382350
rect 331054 382294 331122 382350
rect 331178 382294 361718 382350
rect 361774 382294 361842 382350
rect 361898 382294 392438 382350
rect 392494 382294 392562 382350
rect 392618 382294 423158 382350
rect 423214 382294 423282 382350
rect 423338 382294 453878 382350
rect 453934 382294 454002 382350
rect 454058 382294 484598 382350
rect 484654 382294 484722 382350
rect 484778 382294 515318 382350
rect 515374 382294 515442 382350
rect 515498 382294 546038 382350
rect 546094 382294 546162 382350
rect 546218 382294 561250 382350
rect 561306 382294 561374 382350
rect 561430 382294 561498 382350
rect 561554 382294 561622 382350
rect 561678 382294 579250 382350
rect 579306 382294 579374 382350
rect 579430 382294 579498 382350
rect 579554 382294 579622 382350
rect 579678 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597980 382350
rect -1916 382226 597980 382294
rect -1916 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 3250 382226
rect 3306 382170 3374 382226
rect 3430 382170 3498 382226
rect 3554 382170 3622 382226
rect 3678 382170 21250 382226
rect 21306 382170 21374 382226
rect 21430 382170 21498 382226
rect 21554 382170 21622 382226
rect 21678 382170 39250 382226
rect 39306 382170 39374 382226
rect 39430 382170 39498 382226
rect 39554 382170 39622 382226
rect 39678 382170 54518 382226
rect 54574 382170 54642 382226
rect 54698 382170 57250 382226
rect 57306 382170 57374 382226
rect 57430 382170 57498 382226
rect 57554 382170 57622 382226
rect 57678 382170 75250 382226
rect 75306 382170 75374 382226
rect 75430 382170 75498 382226
rect 75554 382170 75622 382226
rect 75678 382170 85238 382226
rect 85294 382170 85362 382226
rect 85418 382170 93250 382226
rect 93306 382170 93374 382226
rect 93430 382170 93498 382226
rect 93554 382170 93622 382226
rect 93678 382170 111250 382226
rect 111306 382170 111374 382226
rect 111430 382170 111498 382226
rect 111554 382170 111622 382226
rect 111678 382170 115958 382226
rect 116014 382170 116082 382226
rect 116138 382170 146678 382226
rect 146734 382170 146802 382226
rect 146858 382170 177398 382226
rect 177454 382170 177522 382226
rect 177578 382170 208118 382226
rect 208174 382170 208242 382226
rect 208298 382170 238838 382226
rect 238894 382170 238962 382226
rect 239018 382170 269558 382226
rect 269614 382170 269682 382226
rect 269738 382170 300278 382226
rect 300334 382170 300402 382226
rect 300458 382170 330998 382226
rect 331054 382170 331122 382226
rect 331178 382170 361718 382226
rect 361774 382170 361842 382226
rect 361898 382170 392438 382226
rect 392494 382170 392562 382226
rect 392618 382170 423158 382226
rect 423214 382170 423282 382226
rect 423338 382170 453878 382226
rect 453934 382170 454002 382226
rect 454058 382170 484598 382226
rect 484654 382170 484722 382226
rect 484778 382170 515318 382226
rect 515374 382170 515442 382226
rect 515498 382170 546038 382226
rect 546094 382170 546162 382226
rect 546218 382170 561250 382226
rect 561306 382170 561374 382226
rect 561430 382170 561498 382226
rect 561554 382170 561622 382226
rect 561678 382170 579250 382226
rect 579306 382170 579374 382226
rect 579430 382170 579498 382226
rect 579554 382170 579622 382226
rect 579678 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597980 382226
rect -1916 382102 597980 382170
rect -1916 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 3250 382102
rect 3306 382046 3374 382102
rect 3430 382046 3498 382102
rect 3554 382046 3622 382102
rect 3678 382046 21250 382102
rect 21306 382046 21374 382102
rect 21430 382046 21498 382102
rect 21554 382046 21622 382102
rect 21678 382046 39250 382102
rect 39306 382046 39374 382102
rect 39430 382046 39498 382102
rect 39554 382046 39622 382102
rect 39678 382046 54518 382102
rect 54574 382046 54642 382102
rect 54698 382046 57250 382102
rect 57306 382046 57374 382102
rect 57430 382046 57498 382102
rect 57554 382046 57622 382102
rect 57678 382046 75250 382102
rect 75306 382046 75374 382102
rect 75430 382046 75498 382102
rect 75554 382046 75622 382102
rect 75678 382046 85238 382102
rect 85294 382046 85362 382102
rect 85418 382046 93250 382102
rect 93306 382046 93374 382102
rect 93430 382046 93498 382102
rect 93554 382046 93622 382102
rect 93678 382046 111250 382102
rect 111306 382046 111374 382102
rect 111430 382046 111498 382102
rect 111554 382046 111622 382102
rect 111678 382046 115958 382102
rect 116014 382046 116082 382102
rect 116138 382046 146678 382102
rect 146734 382046 146802 382102
rect 146858 382046 177398 382102
rect 177454 382046 177522 382102
rect 177578 382046 208118 382102
rect 208174 382046 208242 382102
rect 208298 382046 238838 382102
rect 238894 382046 238962 382102
rect 239018 382046 269558 382102
rect 269614 382046 269682 382102
rect 269738 382046 300278 382102
rect 300334 382046 300402 382102
rect 300458 382046 330998 382102
rect 331054 382046 331122 382102
rect 331178 382046 361718 382102
rect 361774 382046 361842 382102
rect 361898 382046 392438 382102
rect 392494 382046 392562 382102
rect 392618 382046 423158 382102
rect 423214 382046 423282 382102
rect 423338 382046 453878 382102
rect 453934 382046 454002 382102
rect 454058 382046 484598 382102
rect 484654 382046 484722 382102
rect 484778 382046 515318 382102
rect 515374 382046 515442 382102
rect 515498 382046 546038 382102
rect 546094 382046 546162 382102
rect 546218 382046 561250 382102
rect 561306 382046 561374 382102
rect 561430 382046 561498 382102
rect 561554 382046 561622 382102
rect 561678 382046 579250 382102
rect 579306 382046 579374 382102
rect 579430 382046 579498 382102
rect 579554 382046 579622 382102
rect 579678 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597980 382102
rect -1916 381978 597980 382046
rect -1916 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 3250 381978
rect 3306 381922 3374 381978
rect 3430 381922 3498 381978
rect 3554 381922 3622 381978
rect 3678 381922 21250 381978
rect 21306 381922 21374 381978
rect 21430 381922 21498 381978
rect 21554 381922 21622 381978
rect 21678 381922 39250 381978
rect 39306 381922 39374 381978
rect 39430 381922 39498 381978
rect 39554 381922 39622 381978
rect 39678 381922 54518 381978
rect 54574 381922 54642 381978
rect 54698 381922 57250 381978
rect 57306 381922 57374 381978
rect 57430 381922 57498 381978
rect 57554 381922 57622 381978
rect 57678 381922 75250 381978
rect 75306 381922 75374 381978
rect 75430 381922 75498 381978
rect 75554 381922 75622 381978
rect 75678 381922 85238 381978
rect 85294 381922 85362 381978
rect 85418 381922 93250 381978
rect 93306 381922 93374 381978
rect 93430 381922 93498 381978
rect 93554 381922 93622 381978
rect 93678 381922 111250 381978
rect 111306 381922 111374 381978
rect 111430 381922 111498 381978
rect 111554 381922 111622 381978
rect 111678 381922 115958 381978
rect 116014 381922 116082 381978
rect 116138 381922 146678 381978
rect 146734 381922 146802 381978
rect 146858 381922 177398 381978
rect 177454 381922 177522 381978
rect 177578 381922 208118 381978
rect 208174 381922 208242 381978
rect 208298 381922 238838 381978
rect 238894 381922 238962 381978
rect 239018 381922 269558 381978
rect 269614 381922 269682 381978
rect 269738 381922 300278 381978
rect 300334 381922 300402 381978
rect 300458 381922 330998 381978
rect 331054 381922 331122 381978
rect 331178 381922 361718 381978
rect 361774 381922 361842 381978
rect 361898 381922 392438 381978
rect 392494 381922 392562 381978
rect 392618 381922 423158 381978
rect 423214 381922 423282 381978
rect 423338 381922 453878 381978
rect 453934 381922 454002 381978
rect 454058 381922 484598 381978
rect 484654 381922 484722 381978
rect 484778 381922 515318 381978
rect 515374 381922 515442 381978
rect 515498 381922 546038 381978
rect 546094 381922 546162 381978
rect 546218 381922 561250 381978
rect 561306 381922 561374 381978
rect 561430 381922 561498 381978
rect 561554 381922 561622 381978
rect 561678 381922 579250 381978
rect 579306 381922 579374 381978
rect 579430 381922 579498 381978
rect 579554 381922 579622 381978
rect 579678 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597980 381978
rect -1916 381826 597980 381922
rect -1916 370350 597980 370446
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 6970 370350
rect 7026 370294 7094 370350
rect 7150 370294 7218 370350
rect 7274 370294 7342 370350
rect 7398 370294 24970 370350
rect 25026 370294 25094 370350
rect 25150 370294 25218 370350
rect 25274 370294 25342 370350
rect 25398 370294 42970 370350
rect 43026 370294 43094 370350
rect 43150 370294 43218 370350
rect 43274 370294 43342 370350
rect 43398 370294 60970 370350
rect 61026 370294 61094 370350
rect 61150 370294 61218 370350
rect 61274 370294 61342 370350
rect 61398 370294 69878 370350
rect 69934 370294 70002 370350
rect 70058 370294 78970 370350
rect 79026 370294 79094 370350
rect 79150 370294 79218 370350
rect 79274 370294 79342 370350
rect 79398 370294 96970 370350
rect 97026 370294 97094 370350
rect 97150 370294 97218 370350
rect 97274 370294 97342 370350
rect 97398 370294 100598 370350
rect 100654 370294 100722 370350
rect 100778 370294 131318 370350
rect 131374 370294 131442 370350
rect 131498 370294 162038 370350
rect 162094 370294 162162 370350
rect 162218 370294 192758 370350
rect 192814 370294 192882 370350
rect 192938 370294 223478 370350
rect 223534 370294 223602 370350
rect 223658 370294 254198 370350
rect 254254 370294 254322 370350
rect 254378 370294 284918 370350
rect 284974 370294 285042 370350
rect 285098 370294 315638 370350
rect 315694 370294 315762 370350
rect 315818 370294 346358 370350
rect 346414 370294 346482 370350
rect 346538 370294 377078 370350
rect 377134 370294 377202 370350
rect 377258 370294 407798 370350
rect 407854 370294 407922 370350
rect 407978 370294 438518 370350
rect 438574 370294 438642 370350
rect 438698 370294 469238 370350
rect 469294 370294 469362 370350
rect 469418 370294 499958 370350
rect 500014 370294 500082 370350
rect 500138 370294 530678 370350
rect 530734 370294 530802 370350
rect 530858 370294 564970 370350
rect 565026 370294 565094 370350
rect 565150 370294 565218 370350
rect 565274 370294 565342 370350
rect 565398 370294 582970 370350
rect 583026 370294 583094 370350
rect 583150 370294 583218 370350
rect 583274 370294 583342 370350
rect 583398 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect -1916 370226 597980 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 6970 370226
rect 7026 370170 7094 370226
rect 7150 370170 7218 370226
rect 7274 370170 7342 370226
rect 7398 370170 24970 370226
rect 25026 370170 25094 370226
rect 25150 370170 25218 370226
rect 25274 370170 25342 370226
rect 25398 370170 42970 370226
rect 43026 370170 43094 370226
rect 43150 370170 43218 370226
rect 43274 370170 43342 370226
rect 43398 370170 60970 370226
rect 61026 370170 61094 370226
rect 61150 370170 61218 370226
rect 61274 370170 61342 370226
rect 61398 370170 69878 370226
rect 69934 370170 70002 370226
rect 70058 370170 78970 370226
rect 79026 370170 79094 370226
rect 79150 370170 79218 370226
rect 79274 370170 79342 370226
rect 79398 370170 96970 370226
rect 97026 370170 97094 370226
rect 97150 370170 97218 370226
rect 97274 370170 97342 370226
rect 97398 370170 100598 370226
rect 100654 370170 100722 370226
rect 100778 370170 131318 370226
rect 131374 370170 131442 370226
rect 131498 370170 162038 370226
rect 162094 370170 162162 370226
rect 162218 370170 192758 370226
rect 192814 370170 192882 370226
rect 192938 370170 223478 370226
rect 223534 370170 223602 370226
rect 223658 370170 254198 370226
rect 254254 370170 254322 370226
rect 254378 370170 284918 370226
rect 284974 370170 285042 370226
rect 285098 370170 315638 370226
rect 315694 370170 315762 370226
rect 315818 370170 346358 370226
rect 346414 370170 346482 370226
rect 346538 370170 377078 370226
rect 377134 370170 377202 370226
rect 377258 370170 407798 370226
rect 407854 370170 407922 370226
rect 407978 370170 438518 370226
rect 438574 370170 438642 370226
rect 438698 370170 469238 370226
rect 469294 370170 469362 370226
rect 469418 370170 499958 370226
rect 500014 370170 500082 370226
rect 500138 370170 530678 370226
rect 530734 370170 530802 370226
rect 530858 370170 564970 370226
rect 565026 370170 565094 370226
rect 565150 370170 565218 370226
rect 565274 370170 565342 370226
rect 565398 370170 582970 370226
rect 583026 370170 583094 370226
rect 583150 370170 583218 370226
rect 583274 370170 583342 370226
rect 583398 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect -1916 370102 597980 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 6970 370102
rect 7026 370046 7094 370102
rect 7150 370046 7218 370102
rect 7274 370046 7342 370102
rect 7398 370046 24970 370102
rect 25026 370046 25094 370102
rect 25150 370046 25218 370102
rect 25274 370046 25342 370102
rect 25398 370046 42970 370102
rect 43026 370046 43094 370102
rect 43150 370046 43218 370102
rect 43274 370046 43342 370102
rect 43398 370046 60970 370102
rect 61026 370046 61094 370102
rect 61150 370046 61218 370102
rect 61274 370046 61342 370102
rect 61398 370046 69878 370102
rect 69934 370046 70002 370102
rect 70058 370046 78970 370102
rect 79026 370046 79094 370102
rect 79150 370046 79218 370102
rect 79274 370046 79342 370102
rect 79398 370046 96970 370102
rect 97026 370046 97094 370102
rect 97150 370046 97218 370102
rect 97274 370046 97342 370102
rect 97398 370046 100598 370102
rect 100654 370046 100722 370102
rect 100778 370046 131318 370102
rect 131374 370046 131442 370102
rect 131498 370046 162038 370102
rect 162094 370046 162162 370102
rect 162218 370046 192758 370102
rect 192814 370046 192882 370102
rect 192938 370046 223478 370102
rect 223534 370046 223602 370102
rect 223658 370046 254198 370102
rect 254254 370046 254322 370102
rect 254378 370046 284918 370102
rect 284974 370046 285042 370102
rect 285098 370046 315638 370102
rect 315694 370046 315762 370102
rect 315818 370046 346358 370102
rect 346414 370046 346482 370102
rect 346538 370046 377078 370102
rect 377134 370046 377202 370102
rect 377258 370046 407798 370102
rect 407854 370046 407922 370102
rect 407978 370046 438518 370102
rect 438574 370046 438642 370102
rect 438698 370046 469238 370102
rect 469294 370046 469362 370102
rect 469418 370046 499958 370102
rect 500014 370046 500082 370102
rect 500138 370046 530678 370102
rect 530734 370046 530802 370102
rect 530858 370046 564970 370102
rect 565026 370046 565094 370102
rect 565150 370046 565218 370102
rect 565274 370046 565342 370102
rect 565398 370046 582970 370102
rect 583026 370046 583094 370102
rect 583150 370046 583218 370102
rect 583274 370046 583342 370102
rect 583398 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect -1916 369978 597980 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 6970 369978
rect 7026 369922 7094 369978
rect 7150 369922 7218 369978
rect 7274 369922 7342 369978
rect 7398 369922 24970 369978
rect 25026 369922 25094 369978
rect 25150 369922 25218 369978
rect 25274 369922 25342 369978
rect 25398 369922 42970 369978
rect 43026 369922 43094 369978
rect 43150 369922 43218 369978
rect 43274 369922 43342 369978
rect 43398 369922 60970 369978
rect 61026 369922 61094 369978
rect 61150 369922 61218 369978
rect 61274 369922 61342 369978
rect 61398 369922 69878 369978
rect 69934 369922 70002 369978
rect 70058 369922 78970 369978
rect 79026 369922 79094 369978
rect 79150 369922 79218 369978
rect 79274 369922 79342 369978
rect 79398 369922 96970 369978
rect 97026 369922 97094 369978
rect 97150 369922 97218 369978
rect 97274 369922 97342 369978
rect 97398 369922 100598 369978
rect 100654 369922 100722 369978
rect 100778 369922 131318 369978
rect 131374 369922 131442 369978
rect 131498 369922 162038 369978
rect 162094 369922 162162 369978
rect 162218 369922 192758 369978
rect 192814 369922 192882 369978
rect 192938 369922 223478 369978
rect 223534 369922 223602 369978
rect 223658 369922 254198 369978
rect 254254 369922 254322 369978
rect 254378 369922 284918 369978
rect 284974 369922 285042 369978
rect 285098 369922 315638 369978
rect 315694 369922 315762 369978
rect 315818 369922 346358 369978
rect 346414 369922 346482 369978
rect 346538 369922 377078 369978
rect 377134 369922 377202 369978
rect 377258 369922 407798 369978
rect 407854 369922 407922 369978
rect 407978 369922 438518 369978
rect 438574 369922 438642 369978
rect 438698 369922 469238 369978
rect 469294 369922 469362 369978
rect 469418 369922 499958 369978
rect 500014 369922 500082 369978
rect 500138 369922 530678 369978
rect 530734 369922 530802 369978
rect 530858 369922 564970 369978
rect 565026 369922 565094 369978
rect 565150 369922 565218 369978
rect 565274 369922 565342 369978
rect 565398 369922 582970 369978
rect 583026 369922 583094 369978
rect 583150 369922 583218 369978
rect 583274 369922 583342 369978
rect 583398 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect -1916 369826 597980 369922
rect -1916 364350 597980 364446
rect -1916 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 3250 364350
rect 3306 364294 3374 364350
rect 3430 364294 3498 364350
rect 3554 364294 3622 364350
rect 3678 364294 21250 364350
rect 21306 364294 21374 364350
rect 21430 364294 21498 364350
rect 21554 364294 21622 364350
rect 21678 364294 39250 364350
rect 39306 364294 39374 364350
rect 39430 364294 39498 364350
rect 39554 364294 39622 364350
rect 39678 364294 54518 364350
rect 54574 364294 54642 364350
rect 54698 364294 57250 364350
rect 57306 364294 57374 364350
rect 57430 364294 57498 364350
rect 57554 364294 57622 364350
rect 57678 364294 75250 364350
rect 75306 364294 75374 364350
rect 75430 364294 75498 364350
rect 75554 364294 75622 364350
rect 75678 364294 85238 364350
rect 85294 364294 85362 364350
rect 85418 364294 93250 364350
rect 93306 364294 93374 364350
rect 93430 364294 93498 364350
rect 93554 364294 93622 364350
rect 93678 364294 111250 364350
rect 111306 364294 111374 364350
rect 111430 364294 111498 364350
rect 111554 364294 111622 364350
rect 111678 364294 115958 364350
rect 116014 364294 116082 364350
rect 116138 364294 146678 364350
rect 146734 364294 146802 364350
rect 146858 364294 177398 364350
rect 177454 364294 177522 364350
rect 177578 364294 208118 364350
rect 208174 364294 208242 364350
rect 208298 364294 238838 364350
rect 238894 364294 238962 364350
rect 239018 364294 269558 364350
rect 269614 364294 269682 364350
rect 269738 364294 300278 364350
rect 300334 364294 300402 364350
rect 300458 364294 330998 364350
rect 331054 364294 331122 364350
rect 331178 364294 361718 364350
rect 361774 364294 361842 364350
rect 361898 364294 392438 364350
rect 392494 364294 392562 364350
rect 392618 364294 423158 364350
rect 423214 364294 423282 364350
rect 423338 364294 453878 364350
rect 453934 364294 454002 364350
rect 454058 364294 484598 364350
rect 484654 364294 484722 364350
rect 484778 364294 515318 364350
rect 515374 364294 515442 364350
rect 515498 364294 546038 364350
rect 546094 364294 546162 364350
rect 546218 364294 561250 364350
rect 561306 364294 561374 364350
rect 561430 364294 561498 364350
rect 561554 364294 561622 364350
rect 561678 364294 579250 364350
rect 579306 364294 579374 364350
rect 579430 364294 579498 364350
rect 579554 364294 579622 364350
rect 579678 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597980 364350
rect -1916 364226 597980 364294
rect -1916 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 3250 364226
rect 3306 364170 3374 364226
rect 3430 364170 3498 364226
rect 3554 364170 3622 364226
rect 3678 364170 21250 364226
rect 21306 364170 21374 364226
rect 21430 364170 21498 364226
rect 21554 364170 21622 364226
rect 21678 364170 39250 364226
rect 39306 364170 39374 364226
rect 39430 364170 39498 364226
rect 39554 364170 39622 364226
rect 39678 364170 54518 364226
rect 54574 364170 54642 364226
rect 54698 364170 57250 364226
rect 57306 364170 57374 364226
rect 57430 364170 57498 364226
rect 57554 364170 57622 364226
rect 57678 364170 75250 364226
rect 75306 364170 75374 364226
rect 75430 364170 75498 364226
rect 75554 364170 75622 364226
rect 75678 364170 85238 364226
rect 85294 364170 85362 364226
rect 85418 364170 93250 364226
rect 93306 364170 93374 364226
rect 93430 364170 93498 364226
rect 93554 364170 93622 364226
rect 93678 364170 111250 364226
rect 111306 364170 111374 364226
rect 111430 364170 111498 364226
rect 111554 364170 111622 364226
rect 111678 364170 115958 364226
rect 116014 364170 116082 364226
rect 116138 364170 146678 364226
rect 146734 364170 146802 364226
rect 146858 364170 177398 364226
rect 177454 364170 177522 364226
rect 177578 364170 208118 364226
rect 208174 364170 208242 364226
rect 208298 364170 238838 364226
rect 238894 364170 238962 364226
rect 239018 364170 269558 364226
rect 269614 364170 269682 364226
rect 269738 364170 300278 364226
rect 300334 364170 300402 364226
rect 300458 364170 330998 364226
rect 331054 364170 331122 364226
rect 331178 364170 361718 364226
rect 361774 364170 361842 364226
rect 361898 364170 392438 364226
rect 392494 364170 392562 364226
rect 392618 364170 423158 364226
rect 423214 364170 423282 364226
rect 423338 364170 453878 364226
rect 453934 364170 454002 364226
rect 454058 364170 484598 364226
rect 484654 364170 484722 364226
rect 484778 364170 515318 364226
rect 515374 364170 515442 364226
rect 515498 364170 546038 364226
rect 546094 364170 546162 364226
rect 546218 364170 561250 364226
rect 561306 364170 561374 364226
rect 561430 364170 561498 364226
rect 561554 364170 561622 364226
rect 561678 364170 579250 364226
rect 579306 364170 579374 364226
rect 579430 364170 579498 364226
rect 579554 364170 579622 364226
rect 579678 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597980 364226
rect -1916 364102 597980 364170
rect -1916 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 3250 364102
rect 3306 364046 3374 364102
rect 3430 364046 3498 364102
rect 3554 364046 3622 364102
rect 3678 364046 21250 364102
rect 21306 364046 21374 364102
rect 21430 364046 21498 364102
rect 21554 364046 21622 364102
rect 21678 364046 39250 364102
rect 39306 364046 39374 364102
rect 39430 364046 39498 364102
rect 39554 364046 39622 364102
rect 39678 364046 54518 364102
rect 54574 364046 54642 364102
rect 54698 364046 57250 364102
rect 57306 364046 57374 364102
rect 57430 364046 57498 364102
rect 57554 364046 57622 364102
rect 57678 364046 75250 364102
rect 75306 364046 75374 364102
rect 75430 364046 75498 364102
rect 75554 364046 75622 364102
rect 75678 364046 85238 364102
rect 85294 364046 85362 364102
rect 85418 364046 93250 364102
rect 93306 364046 93374 364102
rect 93430 364046 93498 364102
rect 93554 364046 93622 364102
rect 93678 364046 111250 364102
rect 111306 364046 111374 364102
rect 111430 364046 111498 364102
rect 111554 364046 111622 364102
rect 111678 364046 115958 364102
rect 116014 364046 116082 364102
rect 116138 364046 146678 364102
rect 146734 364046 146802 364102
rect 146858 364046 177398 364102
rect 177454 364046 177522 364102
rect 177578 364046 208118 364102
rect 208174 364046 208242 364102
rect 208298 364046 238838 364102
rect 238894 364046 238962 364102
rect 239018 364046 269558 364102
rect 269614 364046 269682 364102
rect 269738 364046 300278 364102
rect 300334 364046 300402 364102
rect 300458 364046 330998 364102
rect 331054 364046 331122 364102
rect 331178 364046 361718 364102
rect 361774 364046 361842 364102
rect 361898 364046 392438 364102
rect 392494 364046 392562 364102
rect 392618 364046 423158 364102
rect 423214 364046 423282 364102
rect 423338 364046 453878 364102
rect 453934 364046 454002 364102
rect 454058 364046 484598 364102
rect 484654 364046 484722 364102
rect 484778 364046 515318 364102
rect 515374 364046 515442 364102
rect 515498 364046 546038 364102
rect 546094 364046 546162 364102
rect 546218 364046 561250 364102
rect 561306 364046 561374 364102
rect 561430 364046 561498 364102
rect 561554 364046 561622 364102
rect 561678 364046 579250 364102
rect 579306 364046 579374 364102
rect 579430 364046 579498 364102
rect 579554 364046 579622 364102
rect 579678 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597980 364102
rect -1916 363978 597980 364046
rect -1916 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 3250 363978
rect 3306 363922 3374 363978
rect 3430 363922 3498 363978
rect 3554 363922 3622 363978
rect 3678 363922 21250 363978
rect 21306 363922 21374 363978
rect 21430 363922 21498 363978
rect 21554 363922 21622 363978
rect 21678 363922 39250 363978
rect 39306 363922 39374 363978
rect 39430 363922 39498 363978
rect 39554 363922 39622 363978
rect 39678 363922 54518 363978
rect 54574 363922 54642 363978
rect 54698 363922 57250 363978
rect 57306 363922 57374 363978
rect 57430 363922 57498 363978
rect 57554 363922 57622 363978
rect 57678 363922 75250 363978
rect 75306 363922 75374 363978
rect 75430 363922 75498 363978
rect 75554 363922 75622 363978
rect 75678 363922 85238 363978
rect 85294 363922 85362 363978
rect 85418 363922 93250 363978
rect 93306 363922 93374 363978
rect 93430 363922 93498 363978
rect 93554 363922 93622 363978
rect 93678 363922 111250 363978
rect 111306 363922 111374 363978
rect 111430 363922 111498 363978
rect 111554 363922 111622 363978
rect 111678 363922 115958 363978
rect 116014 363922 116082 363978
rect 116138 363922 146678 363978
rect 146734 363922 146802 363978
rect 146858 363922 177398 363978
rect 177454 363922 177522 363978
rect 177578 363922 208118 363978
rect 208174 363922 208242 363978
rect 208298 363922 238838 363978
rect 238894 363922 238962 363978
rect 239018 363922 269558 363978
rect 269614 363922 269682 363978
rect 269738 363922 300278 363978
rect 300334 363922 300402 363978
rect 300458 363922 330998 363978
rect 331054 363922 331122 363978
rect 331178 363922 361718 363978
rect 361774 363922 361842 363978
rect 361898 363922 392438 363978
rect 392494 363922 392562 363978
rect 392618 363922 423158 363978
rect 423214 363922 423282 363978
rect 423338 363922 453878 363978
rect 453934 363922 454002 363978
rect 454058 363922 484598 363978
rect 484654 363922 484722 363978
rect 484778 363922 515318 363978
rect 515374 363922 515442 363978
rect 515498 363922 546038 363978
rect 546094 363922 546162 363978
rect 546218 363922 561250 363978
rect 561306 363922 561374 363978
rect 561430 363922 561498 363978
rect 561554 363922 561622 363978
rect 561678 363922 579250 363978
rect 579306 363922 579374 363978
rect 579430 363922 579498 363978
rect 579554 363922 579622 363978
rect 579678 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597980 363978
rect -1916 363826 597980 363922
rect -1916 352350 597980 352446
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 6970 352350
rect 7026 352294 7094 352350
rect 7150 352294 7218 352350
rect 7274 352294 7342 352350
rect 7398 352294 24970 352350
rect 25026 352294 25094 352350
rect 25150 352294 25218 352350
rect 25274 352294 25342 352350
rect 25398 352294 42970 352350
rect 43026 352294 43094 352350
rect 43150 352294 43218 352350
rect 43274 352294 43342 352350
rect 43398 352294 60970 352350
rect 61026 352294 61094 352350
rect 61150 352294 61218 352350
rect 61274 352294 61342 352350
rect 61398 352294 69878 352350
rect 69934 352294 70002 352350
rect 70058 352294 78970 352350
rect 79026 352294 79094 352350
rect 79150 352294 79218 352350
rect 79274 352294 79342 352350
rect 79398 352294 96970 352350
rect 97026 352294 97094 352350
rect 97150 352294 97218 352350
rect 97274 352294 97342 352350
rect 97398 352294 100598 352350
rect 100654 352294 100722 352350
rect 100778 352294 131318 352350
rect 131374 352294 131442 352350
rect 131498 352294 162038 352350
rect 162094 352294 162162 352350
rect 162218 352294 192758 352350
rect 192814 352294 192882 352350
rect 192938 352294 223478 352350
rect 223534 352294 223602 352350
rect 223658 352294 254198 352350
rect 254254 352294 254322 352350
rect 254378 352294 284918 352350
rect 284974 352294 285042 352350
rect 285098 352294 315638 352350
rect 315694 352294 315762 352350
rect 315818 352294 346358 352350
rect 346414 352294 346482 352350
rect 346538 352294 377078 352350
rect 377134 352294 377202 352350
rect 377258 352294 407798 352350
rect 407854 352294 407922 352350
rect 407978 352294 438518 352350
rect 438574 352294 438642 352350
rect 438698 352294 469238 352350
rect 469294 352294 469362 352350
rect 469418 352294 499958 352350
rect 500014 352294 500082 352350
rect 500138 352294 530678 352350
rect 530734 352294 530802 352350
rect 530858 352294 564970 352350
rect 565026 352294 565094 352350
rect 565150 352294 565218 352350
rect 565274 352294 565342 352350
rect 565398 352294 582970 352350
rect 583026 352294 583094 352350
rect 583150 352294 583218 352350
rect 583274 352294 583342 352350
rect 583398 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect -1916 352226 597980 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 6970 352226
rect 7026 352170 7094 352226
rect 7150 352170 7218 352226
rect 7274 352170 7342 352226
rect 7398 352170 24970 352226
rect 25026 352170 25094 352226
rect 25150 352170 25218 352226
rect 25274 352170 25342 352226
rect 25398 352170 42970 352226
rect 43026 352170 43094 352226
rect 43150 352170 43218 352226
rect 43274 352170 43342 352226
rect 43398 352170 60970 352226
rect 61026 352170 61094 352226
rect 61150 352170 61218 352226
rect 61274 352170 61342 352226
rect 61398 352170 69878 352226
rect 69934 352170 70002 352226
rect 70058 352170 78970 352226
rect 79026 352170 79094 352226
rect 79150 352170 79218 352226
rect 79274 352170 79342 352226
rect 79398 352170 96970 352226
rect 97026 352170 97094 352226
rect 97150 352170 97218 352226
rect 97274 352170 97342 352226
rect 97398 352170 100598 352226
rect 100654 352170 100722 352226
rect 100778 352170 131318 352226
rect 131374 352170 131442 352226
rect 131498 352170 162038 352226
rect 162094 352170 162162 352226
rect 162218 352170 192758 352226
rect 192814 352170 192882 352226
rect 192938 352170 223478 352226
rect 223534 352170 223602 352226
rect 223658 352170 254198 352226
rect 254254 352170 254322 352226
rect 254378 352170 284918 352226
rect 284974 352170 285042 352226
rect 285098 352170 315638 352226
rect 315694 352170 315762 352226
rect 315818 352170 346358 352226
rect 346414 352170 346482 352226
rect 346538 352170 377078 352226
rect 377134 352170 377202 352226
rect 377258 352170 407798 352226
rect 407854 352170 407922 352226
rect 407978 352170 438518 352226
rect 438574 352170 438642 352226
rect 438698 352170 469238 352226
rect 469294 352170 469362 352226
rect 469418 352170 499958 352226
rect 500014 352170 500082 352226
rect 500138 352170 530678 352226
rect 530734 352170 530802 352226
rect 530858 352170 564970 352226
rect 565026 352170 565094 352226
rect 565150 352170 565218 352226
rect 565274 352170 565342 352226
rect 565398 352170 582970 352226
rect 583026 352170 583094 352226
rect 583150 352170 583218 352226
rect 583274 352170 583342 352226
rect 583398 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect -1916 352102 597980 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 6970 352102
rect 7026 352046 7094 352102
rect 7150 352046 7218 352102
rect 7274 352046 7342 352102
rect 7398 352046 24970 352102
rect 25026 352046 25094 352102
rect 25150 352046 25218 352102
rect 25274 352046 25342 352102
rect 25398 352046 42970 352102
rect 43026 352046 43094 352102
rect 43150 352046 43218 352102
rect 43274 352046 43342 352102
rect 43398 352046 60970 352102
rect 61026 352046 61094 352102
rect 61150 352046 61218 352102
rect 61274 352046 61342 352102
rect 61398 352046 69878 352102
rect 69934 352046 70002 352102
rect 70058 352046 78970 352102
rect 79026 352046 79094 352102
rect 79150 352046 79218 352102
rect 79274 352046 79342 352102
rect 79398 352046 96970 352102
rect 97026 352046 97094 352102
rect 97150 352046 97218 352102
rect 97274 352046 97342 352102
rect 97398 352046 100598 352102
rect 100654 352046 100722 352102
rect 100778 352046 131318 352102
rect 131374 352046 131442 352102
rect 131498 352046 162038 352102
rect 162094 352046 162162 352102
rect 162218 352046 192758 352102
rect 192814 352046 192882 352102
rect 192938 352046 223478 352102
rect 223534 352046 223602 352102
rect 223658 352046 254198 352102
rect 254254 352046 254322 352102
rect 254378 352046 284918 352102
rect 284974 352046 285042 352102
rect 285098 352046 315638 352102
rect 315694 352046 315762 352102
rect 315818 352046 346358 352102
rect 346414 352046 346482 352102
rect 346538 352046 377078 352102
rect 377134 352046 377202 352102
rect 377258 352046 407798 352102
rect 407854 352046 407922 352102
rect 407978 352046 438518 352102
rect 438574 352046 438642 352102
rect 438698 352046 469238 352102
rect 469294 352046 469362 352102
rect 469418 352046 499958 352102
rect 500014 352046 500082 352102
rect 500138 352046 530678 352102
rect 530734 352046 530802 352102
rect 530858 352046 564970 352102
rect 565026 352046 565094 352102
rect 565150 352046 565218 352102
rect 565274 352046 565342 352102
rect 565398 352046 582970 352102
rect 583026 352046 583094 352102
rect 583150 352046 583218 352102
rect 583274 352046 583342 352102
rect 583398 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect -1916 351978 597980 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 6970 351978
rect 7026 351922 7094 351978
rect 7150 351922 7218 351978
rect 7274 351922 7342 351978
rect 7398 351922 24970 351978
rect 25026 351922 25094 351978
rect 25150 351922 25218 351978
rect 25274 351922 25342 351978
rect 25398 351922 42970 351978
rect 43026 351922 43094 351978
rect 43150 351922 43218 351978
rect 43274 351922 43342 351978
rect 43398 351922 60970 351978
rect 61026 351922 61094 351978
rect 61150 351922 61218 351978
rect 61274 351922 61342 351978
rect 61398 351922 69878 351978
rect 69934 351922 70002 351978
rect 70058 351922 78970 351978
rect 79026 351922 79094 351978
rect 79150 351922 79218 351978
rect 79274 351922 79342 351978
rect 79398 351922 96970 351978
rect 97026 351922 97094 351978
rect 97150 351922 97218 351978
rect 97274 351922 97342 351978
rect 97398 351922 100598 351978
rect 100654 351922 100722 351978
rect 100778 351922 131318 351978
rect 131374 351922 131442 351978
rect 131498 351922 162038 351978
rect 162094 351922 162162 351978
rect 162218 351922 192758 351978
rect 192814 351922 192882 351978
rect 192938 351922 223478 351978
rect 223534 351922 223602 351978
rect 223658 351922 254198 351978
rect 254254 351922 254322 351978
rect 254378 351922 284918 351978
rect 284974 351922 285042 351978
rect 285098 351922 315638 351978
rect 315694 351922 315762 351978
rect 315818 351922 346358 351978
rect 346414 351922 346482 351978
rect 346538 351922 377078 351978
rect 377134 351922 377202 351978
rect 377258 351922 407798 351978
rect 407854 351922 407922 351978
rect 407978 351922 438518 351978
rect 438574 351922 438642 351978
rect 438698 351922 469238 351978
rect 469294 351922 469362 351978
rect 469418 351922 499958 351978
rect 500014 351922 500082 351978
rect 500138 351922 530678 351978
rect 530734 351922 530802 351978
rect 530858 351922 564970 351978
rect 565026 351922 565094 351978
rect 565150 351922 565218 351978
rect 565274 351922 565342 351978
rect 565398 351922 582970 351978
rect 583026 351922 583094 351978
rect 583150 351922 583218 351978
rect 583274 351922 583342 351978
rect 583398 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect -1916 351826 597980 351922
rect -1916 346350 597980 346446
rect -1916 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 3250 346350
rect 3306 346294 3374 346350
rect 3430 346294 3498 346350
rect 3554 346294 3622 346350
rect 3678 346294 21250 346350
rect 21306 346294 21374 346350
rect 21430 346294 21498 346350
rect 21554 346294 21622 346350
rect 21678 346294 39250 346350
rect 39306 346294 39374 346350
rect 39430 346294 39498 346350
rect 39554 346294 39622 346350
rect 39678 346294 54518 346350
rect 54574 346294 54642 346350
rect 54698 346294 57250 346350
rect 57306 346294 57374 346350
rect 57430 346294 57498 346350
rect 57554 346294 57622 346350
rect 57678 346294 75250 346350
rect 75306 346294 75374 346350
rect 75430 346294 75498 346350
rect 75554 346294 75622 346350
rect 75678 346294 85238 346350
rect 85294 346294 85362 346350
rect 85418 346294 93250 346350
rect 93306 346294 93374 346350
rect 93430 346294 93498 346350
rect 93554 346294 93622 346350
rect 93678 346294 111250 346350
rect 111306 346294 111374 346350
rect 111430 346294 111498 346350
rect 111554 346294 111622 346350
rect 111678 346294 115958 346350
rect 116014 346294 116082 346350
rect 116138 346294 146678 346350
rect 146734 346294 146802 346350
rect 146858 346294 177398 346350
rect 177454 346294 177522 346350
rect 177578 346294 208118 346350
rect 208174 346294 208242 346350
rect 208298 346294 238838 346350
rect 238894 346294 238962 346350
rect 239018 346294 269558 346350
rect 269614 346294 269682 346350
rect 269738 346294 300278 346350
rect 300334 346294 300402 346350
rect 300458 346294 330998 346350
rect 331054 346294 331122 346350
rect 331178 346294 361718 346350
rect 361774 346294 361842 346350
rect 361898 346294 392438 346350
rect 392494 346294 392562 346350
rect 392618 346294 423158 346350
rect 423214 346294 423282 346350
rect 423338 346294 453878 346350
rect 453934 346294 454002 346350
rect 454058 346294 484598 346350
rect 484654 346294 484722 346350
rect 484778 346294 515318 346350
rect 515374 346294 515442 346350
rect 515498 346294 546038 346350
rect 546094 346294 546162 346350
rect 546218 346294 561250 346350
rect 561306 346294 561374 346350
rect 561430 346294 561498 346350
rect 561554 346294 561622 346350
rect 561678 346294 579250 346350
rect 579306 346294 579374 346350
rect 579430 346294 579498 346350
rect 579554 346294 579622 346350
rect 579678 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597980 346350
rect -1916 346226 597980 346294
rect -1916 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 3250 346226
rect 3306 346170 3374 346226
rect 3430 346170 3498 346226
rect 3554 346170 3622 346226
rect 3678 346170 21250 346226
rect 21306 346170 21374 346226
rect 21430 346170 21498 346226
rect 21554 346170 21622 346226
rect 21678 346170 39250 346226
rect 39306 346170 39374 346226
rect 39430 346170 39498 346226
rect 39554 346170 39622 346226
rect 39678 346170 54518 346226
rect 54574 346170 54642 346226
rect 54698 346170 57250 346226
rect 57306 346170 57374 346226
rect 57430 346170 57498 346226
rect 57554 346170 57622 346226
rect 57678 346170 75250 346226
rect 75306 346170 75374 346226
rect 75430 346170 75498 346226
rect 75554 346170 75622 346226
rect 75678 346170 85238 346226
rect 85294 346170 85362 346226
rect 85418 346170 93250 346226
rect 93306 346170 93374 346226
rect 93430 346170 93498 346226
rect 93554 346170 93622 346226
rect 93678 346170 111250 346226
rect 111306 346170 111374 346226
rect 111430 346170 111498 346226
rect 111554 346170 111622 346226
rect 111678 346170 115958 346226
rect 116014 346170 116082 346226
rect 116138 346170 146678 346226
rect 146734 346170 146802 346226
rect 146858 346170 177398 346226
rect 177454 346170 177522 346226
rect 177578 346170 208118 346226
rect 208174 346170 208242 346226
rect 208298 346170 238838 346226
rect 238894 346170 238962 346226
rect 239018 346170 269558 346226
rect 269614 346170 269682 346226
rect 269738 346170 300278 346226
rect 300334 346170 300402 346226
rect 300458 346170 330998 346226
rect 331054 346170 331122 346226
rect 331178 346170 361718 346226
rect 361774 346170 361842 346226
rect 361898 346170 392438 346226
rect 392494 346170 392562 346226
rect 392618 346170 423158 346226
rect 423214 346170 423282 346226
rect 423338 346170 453878 346226
rect 453934 346170 454002 346226
rect 454058 346170 484598 346226
rect 484654 346170 484722 346226
rect 484778 346170 515318 346226
rect 515374 346170 515442 346226
rect 515498 346170 546038 346226
rect 546094 346170 546162 346226
rect 546218 346170 561250 346226
rect 561306 346170 561374 346226
rect 561430 346170 561498 346226
rect 561554 346170 561622 346226
rect 561678 346170 579250 346226
rect 579306 346170 579374 346226
rect 579430 346170 579498 346226
rect 579554 346170 579622 346226
rect 579678 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597980 346226
rect -1916 346102 597980 346170
rect -1916 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 3250 346102
rect 3306 346046 3374 346102
rect 3430 346046 3498 346102
rect 3554 346046 3622 346102
rect 3678 346046 21250 346102
rect 21306 346046 21374 346102
rect 21430 346046 21498 346102
rect 21554 346046 21622 346102
rect 21678 346046 39250 346102
rect 39306 346046 39374 346102
rect 39430 346046 39498 346102
rect 39554 346046 39622 346102
rect 39678 346046 54518 346102
rect 54574 346046 54642 346102
rect 54698 346046 57250 346102
rect 57306 346046 57374 346102
rect 57430 346046 57498 346102
rect 57554 346046 57622 346102
rect 57678 346046 75250 346102
rect 75306 346046 75374 346102
rect 75430 346046 75498 346102
rect 75554 346046 75622 346102
rect 75678 346046 85238 346102
rect 85294 346046 85362 346102
rect 85418 346046 93250 346102
rect 93306 346046 93374 346102
rect 93430 346046 93498 346102
rect 93554 346046 93622 346102
rect 93678 346046 111250 346102
rect 111306 346046 111374 346102
rect 111430 346046 111498 346102
rect 111554 346046 111622 346102
rect 111678 346046 115958 346102
rect 116014 346046 116082 346102
rect 116138 346046 146678 346102
rect 146734 346046 146802 346102
rect 146858 346046 177398 346102
rect 177454 346046 177522 346102
rect 177578 346046 208118 346102
rect 208174 346046 208242 346102
rect 208298 346046 238838 346102
rect 238894 346046 238962 346102
rect 239018 346046 269558 346102
rect 269614 346046 269682 346102
rect 269738 346046 300278 346102
rect 300334 346046 300402 346102
rect 300458 346046 330998 346102
rect 331054 346046 331122 346102
rect 331178 346046 361718 346102
rect 361774 346046 361842 346102
rect 361898 346046 392438 346102
rect 392494 346046 392562 346102
rect 392618 346046 423158 346102
rect 423214 346046 423282 346102
rect 423338 346046 453878 346102
rect 453934 346046 454002 346102
rect 454058 346046 484598 346102
rect 484654 346046 484722 346102
rect 484778 346046 515318 346102
rect 515374 346046 515442 346102
rect 515498 346046 546038 346102
rect 546094 346046 546162 346102
rect 546218 346046 561250 346102
rect 561306 346046 561374 346102
rect 561430 346046 561498 346102
rect 561554 346046 561622 346102
rect 561678 346046 579250 346102
rect 579306 346046 579374 346102
rect 579430 346046 579498 346102
rect 579554 346046 579622 346102
rect 579678 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597980 346102
rect -1916 345978 597980 346046
rect -1916 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 3250 345978
rect 3306 345922 3374 345978
rect 3430 345922 3498 345978
rect 3554 345922 3622 345978
rect 3678 345922 21250 345978
rect 21306 345922 21374 345978
rect 21430 345922 21498 345978
rect 21554 345922 21622 345978
rect 21678 345922 39250 345978
rect 39306 345922 39374 345978
rect 39430 345922 39498 345978
rect 39554 345922 39622 345978
rect 39678 345922 54518 345978
rect 54574 345922 54642 345978
rect 54698 345922 57250 345978
rect 57306 345922 57374 345978
rect 57430 345922 57498 345978
rect 57554 345922 57622 345978
rect 57678 345922 75250 345978
rect 75306 345922 75374 345978
rect 75430 345922 75498 345978
rect 75554 345922 75622 345978
rect 75678 345922 85238 345978
rect 85294 345922 85362 345978
rect 85418 345922 93250 345978
rect 93306 345922 93374 345978
rect 93430 345922 93498 345978
rect 93554 345922 93622 345978
rect 93678 345922 111250 345978
rect 111306 345922 111374 345978
rect 111430 345922 111498 345978
rect 111554 345922 111622 345978
rect 111678 345922 115958 345978
rect 116014 345922 116082 345978
rect 116138 345922 146678 345978
rect 146734 345922 146802 345978
rect 146858 345922 177398 345978
rect 177454 345922 177522 345978
rect 177578 345922 208118 345978
rect 208174 345922 208242 345978
rect 208298 345922 238838 345978
rect 238894 345922 238962 345978
rect 239018 345922 269558 345978
rect 269614 345922 269682 345978
rect 269738 345922 300278 345978
rect 300334 345922 300402 345978
rect 300458 345922 330998 345978
rect 331054 345922 331122 345978
rect 331178 345922 361718 345978
rect 361774 345922 361842 345978
rect 361898 345922 392438 345978
rect 392494 345922 392562 345978
rect 392618 345922 423158 345978
rect 423214 345922 423282 345978
rect 423338 345922 453878 345978
rect 453934 345922 454002 345978
rect 454058 345922 484598 345978
rect 484654 345922 484722 345978
rect 484778 345922 515318 345978
rect 515374 345922 515442 345978
rect 515498 345922 546038 345978
rect 546094 345922 546162 345978
rect 546218 345922 561250 345978
rect 561306 345922 561374 345978
rect 561430 345922 561498 345978
rect 561554 345922 561622 345978
rect 561678 345922 579250 345978
rect 579306 345922 579374 345978
rect 579430 345922 579498 345978
rect 579554 345922 579622 345978
rect 579678 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597980 345978
rect -1916 345826 597980 345922
rect -1916 334350 597980 334446
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 6970 334350
rect 7026 334294 7094 334350
rect 7150 334294 7218 334350
rect 7274 334294 7342 334350
rect 7398 334294 24970 334350
rect 25026 334294 25094 334350
rect 25150 334294 25218 334350
rect 25274 334294 25342 334350
rect 25398 334294 42970 334350
rect 43026 334294 43094 334350
rect 43150 334294 43218 334350
rect 43274 334294 43342 334350
rect 43398 334294 60970 334350
rect 61026 334294 61094 334350
rect 61150 334294 61218 334350
rect 61274 334294 61342 334350
rect 61398 334294 69878 334350
rect 69934 334294 70002 334350
rect 70058 334294 78970 334350
rect 79026 334294 79094 334350
rect 79150 334294 79218 334350
rect 79274 334294 79342 334350
rect 79398 334294 96970 334350
rect 97026 334294 97094 334350
rect 97150 334294 97218 334350
rect 97274 334294 97342 334350
rect 97398 334294 100598 334350
rect 100654 334294 100722 334350
rect 100778 334294 131318 334350
rect 131374 334294 131442 334350
rect 131498 334294 162038 334350
rect 162094 334294 162162 334350
rect 162218 334294 192758 334350
rect 192814 334294 192882 334350
rect 192938 334294 223478 334350
rect 223534 334294 223602 334350
rect 223658 334294 254198 334350
rect 254254 334294 254322 334350
rect 254378 334294 284918 334350
rect 284974 334294 285042 334350
rect 285098 334294 315638 334350
rect 315694 334294 315762 334350
rect 315818 334294 346358 334350
rect 346414 334294 346482 334350
rect 346538 334294 377078 334350
rect 377134 334294 377202 334350
rect 377258 334294 407798 334350
rect 407854 334294 407922 334350
rect 407978 334294 438518 334350
rect 438574 334294 438642 334350
rect 438698 334294 469238 334350
rect 469294 334294 469362 334350
rect 469418 334294 499958 334350
rect 500014 334294 500082 334350
rect 500138 334294 530678 334350
rect 530734 334294 530802 334350
rect 530858 334294 564970 334350
rect 565026 334294 565094 334350
rect 565150 334294 565218 334350
rect 565274 334294 565342 334350
rect 565398 334294 582970 334350
rect 583026 334294 583094 334350
rect 583150 334294 583218 334350
rect 583274 334294 583342 334350
rect 583398 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect -1916 334226 597980 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 6970 334226
rect 7026 334170 7094 334226
rect 7150 334170 7218 334226
rect 7274 334170 7342 334226
rect 7398 334170 24970 334226
rect 25026 334170 25094 334226
rect 25150 334170 25218 334226
rect 25274 334170 25342 334226
rect 25398 334170 42970 334226
rect 43026 334170 43094 334226
rect 43150 334170 43218 334226
rect 43274 334170 43342 334226
rect 43398 334170 60970 334226
rect 61026 334170 61094 334226
rect 61150 334170 61218 334226
rect 61274 334170 61342 334226
rect 61398 334170 69878 334226
rect 69934 334170 70002 334226
rect 70058 334170 78970 334226
rect 79026 334170 79094 334226
rect 79150 334170 79218 334226
rect 79274 334170 79342 334226
rect 79398 334170 96970 334226
rect 97026 334170 97094 334226
rect 97150 334170 97218 334226
rect 97274 334170 97342 334226
rect 97398 334170 100598 334226
rect 100654 334170 100722 334226
rect 100778 334170 131318 334226
rect 131374 334170 131442 334226
rect 131498 334170 162038 334226
rect 162094 334170 162162 334226
rect 162218 334170 192758 334226
rect 192814 334170 192882 334226
rect 192938 334170 223478 334226
rect 223534 334170 223602 334226
rect 223658 334170 254198 334226
rect 254254 334170 254322 334226
rect 254378 334170 284918 334226
rect 284974 334170 285042 334226
rect 285098 334170 315638 334226
rect 315694 334170 315762 334226
rect 315818 334170 346358 334226
rect 346414 334170 346482 334226
rect 346538 334170 377078 334226
rect 377134 334170 377202 334226
rect 377258 334170 407798 334226
rect 407854 334170 407922 334226
rect 407978 334170 438518 334226
rect 438574 334170 438642 334226
rect 438698 334170 469238 334226
rect 469294 334170 469362 334226
rect 469418 334170 499958 334226
rect 500014 334170 500082 334226
rect 500138 334170 530678 334226
rect 530734 334170 530802 334226
rect 530858 334170 564970 334226
rect 565026 334170 565094 334226
rect 565150 334170 565218 334226
rect 565274 334170 565342 334226
rect 565398 334170 582970 334226
rect 583026 334170 583094 334226
rect 583150 334170 583218 334226
rect 583274 334170 583342 334226
rect 583398 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect -1916 334102 597980 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 6970 334102
rect 7026 334046 7094 334102
rect 7150 334046 7218 334102
rect 7274 334046 7342 334102
rect 7398 334046 24970 334102
rect 25026 334046 25094 334102
rect 25150 334046 25218 334102
rect 25274 334046 25342 334102
rect 25398 334046 42970 334102
rect 43026 334046 43094 334102
rect 43150 334046 43218 334102
rect 43274 334046 43342 334102
rect 43398 334046 60970 334102
rect 61026 334046 61094 334102
rect 61150 334046 61218 334102
rect 61274 334046 61342 334102
rect 61398 334046 69878 334102
rect 69934 334046 70002 334102
rect 70058 334046 78970 334102
rect 79026 334046 79094 334102
rect 79150 334046 79218 334102
rect 79274 334046 79342 334102
rect 79398 334046 96970 334102
rect 97026 334046 97094 334102
rect 97150 334046 97218 334102
rect 97274 334046 97342 334102
rect 97398 334046 100598 334102
rect 100654 334046 100722 334102
rect 100778 334046 131318 334102
rect 131374 334046 131442 334102
rect 131498 334046 162038 334102
rect 162094 334046 162162 334102
rect 162218 334046 192758 334102
rect 192814 334046 192882 334102
rect 192938 334046 223478 334102
rect 223534 334046 223602 334102
rect 223658 334046 254198 334102
rect 254254 334046 254322 334102
rect 254378 334046 284918 334102
rect 284974 334046 285042 334102
rect 285098 334046 315638 334102
rect 315694 334046 315762 334102
rect 315818 334046 346358 334102
rect 346414 334046 346482 334102
rect 346538 334046 377078 334102
rect 377134 334046 377202 334102
rect 377258 334046 407798 334102
rect 407854 334046 407922 334102
rect 407978 334046 438518 334102
rect 438574 334046 438642 334102
rect 438698 334046 469238 334102
rect 469294 334046 469362 334102
rect 469418 334046 499958 334102
rect 500014 334046 500082 334102
rect 500138 334046 530678 334102
rect 530734 334046 530802 334102
rect 530858 334046 564970 334102
rect 565026 334046 565094 334102
rect 565150 334046 565218 334102
rect 565274 334046 565342 334102
rect 565398 334046 582970 334102
rect 583026 334046 583094 334102
rect 583150 334046 583218 334102
rect 583274 334046 583342 334102
rect 583398 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect -1916 333978 597980 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 6970 333978
rect 7026 333922 7094 333978
rect 7150 333922 7218 333978
rect 7274 333922 7342 333978
rect 7398 333922 24970 333978
rect 25026 333922 25094 333978
rect 25150 333922 25218 333978
rect 25274 333922 25342 333978
rect 25398 333922 42970 333978
rect 43026 333922 43094 333978
rect 43150 333922 43218 333978
rect 43274 333922 43342 333978
rect 43398 333922 60970 333978
rect 61026 333922 61094 333978
rect 61150 333922 61218 333978
rect 61274 333922 61342 333978
rect 61398 333922 69878 333978
rect 69934 333922 70002 333978
rect 70058 333922 78970 333978
rect 79026 333922 79094 333978
rect 79150 333922 79218 333978
rect 79274 333922 79342 333978
rect 79398 333922 96970 333978
rect 97026 333922 97094 333978
rect 97150 333922 97218 333978
rect 97274 333922 97342 333978
rect 97398 333922 100598 333978
rect 100654 333922 100722 333978
rect 100778 333922 131318 333978
rect 131374 333922 131442 333978
rect 131498 333922 162038 333978
rect 162094 333922 162162 333978
rect 162218 333922 192758 333978
rect 192814 333922 192882 333978
rect 192938 333922 223478 333978
rect 223534 333922 223602 333978
rect 223658 333922 254198 333978
rect 254254 333922 254322 333978
rect 254378 333922 284918 333978
rect 284974 333922 285042 333978
rect 285098 333922 315638 333978
rect 315694 333922 315762 333978
rect 315818 333922 346358 333978
rect 346414 333922 346482 333978
rect 346538 333922 377078 333978
rect 377134 333922 377202 333978
rect 377258 333922 407798 333978
rect 407854 333922 407922 333978
rect 407978 333922 438518 333978
rect 438574 333922 438642 333978
rect 438698 333922 469238 333978
rect 469294 333922 469362 333978
rect 469418 333922 499958 333978
rect 500014 333922 500082 333978
rect 500138 333922 530678 333978
rect 530734 333922 530802 333978
rect 530858 333922 564970 333978
rect 565026 333922 565094 333978
rect 565150 333922 565218 333978
rect 565274 333922 565342 333978
rect 565398 333922 582970 333978
rect 583026 333922 583094 333978
rect 583150 333922 583218 333978
rect 583274 333922 583342 333978
rect 583398 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect -1916 333826 597980 333922
rect -1916 328350 597980 328446
rect -1916 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 3250 328350
rect 3306 328294 3374 328350
rect 3430 328294 3498 328350
rect 3554 328294 3622 328350
rect 3678 328294 21250 328350
rect 21306 328294 21374 328350
rect 21430 328294 21498 328350
rect 21554 328294 21622 328350
rect 21678 328294 39250 328350
rect 39306 328294 39374 328350
rect 39430 328294 39498 328350
rect 39554 328294 39622 328350
rect 39678 328294 54518 328350
rect 54574 328294 54642 328350
rect 54698 328294 57250 328350
rect 57306 328294 57374 328350
rect 57430 328294 57498 328350
rect 57554 328294 57622 328350
rect 57678 328294 75250 328350
rect 75306 328294 75374 328350
rect 75430 328294 75498 328350
rect 75554 328294 75622 328350
rect 75678 328294 85238 328350
rect 85294 328294 85362 328350
rect 85418 328294 93250 328350
rect 93306 328294 93374 328350
rect 93430 328294 93498 328350
rect 93554 328294 93622 328350
rect 93678 328294 111250 328350
rect 111306 328294 111374 328350
rect 111430 328294 111498 328350
rect 111554 328294 111622 328350
rect 111678 328294 115958 328350
rect 116014 328294 116082 328350
rect 116138 328294 146678 328350
rect 146734 328294 146802 328350
rect 146858 328294 177398 328350
rect 177454 328294 177522 328350
rect 177578 328294 208118 328350
rect 208174 328294 208242 328350
rect 208298 328294 238838 328350
rect 238894 328294 238962 328350
rect 239018 328294 269558 328350
rect 269614 328294 269682 328350
rect 269738 328294 300278 328350
rect 300334 328294 300402 328350
rect 300458 328294 330998 328350
rect 331054 328294 331122 328350
rect 331178 328294 361718 328350
rect 361774 328294 361842 328350
rect 361898 328294 392438 328350
rect 392494 328294 392562 328350
rect 392618 328294 423158 328350
rect 423214 328294 423282 328350
rect 423338 328294 453878 328350
rect 453934 328294 454002 328350
rect 454058 328294 484598 328350
rect 484654 328294 484722 328350
rect 484778 328294 515318 328350
rect 515374 328294 515442 328350
rect 515498 328294 546038 328350
rect 546094 328294 546162 328350
rect 546218 328294 561250 328350
rect 561306 328294 561374 328350
rect 561430 328294 561498 328350
rect 561554 328294 561622 328350
rect 561678 328294 579250 328350
rect 579306 328294 579374 328350
rect 579430 328294 579498 328350
rect 579554 328294 579622 328350
rect 579678 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597980 328350
rect -1916 328226 597980 328294
rect -1916 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 3250 328226
rect 3306 328170 3374 328226
rect 3430 328170 3498 328226
rect 3554 328170 3622 328226
rect 3678 328170 21250 328226
rect 21306 328170 21374 328226
rect 21430 328170 21498 328226
rect 21554 328170 21622 328226
rect 21678 328170 39250 328226
rect 39306 328170 39374 328226
rect 39430 328170 39498 328226
rect 39554 328170 39622 328226
rect 39678 328170 54518 328226
rect 54574 328170 54642 328226
rect 54698 328170 57250 328226
rect 57306 328170 57374 328226
rect 57430 328170 57498 328226
rect 57554 328170 57622 328226
rect 57678 328170 75250 328226
rect 75306 328170 75374 328226
rect 75430 328170 75498 328226
rect 75554 328170 75622 328226
rect 75678 328170 85238 328226
rect 85294 328170 85362 328226
rect 85418 328170 93250 328226
rect 93306 328170 93374 328226
rect 93430 328170 93498 328226
rect 93554 328170 93622 328226
rect 93678 328170 111250 328226
rect 111306 328170 111374 328226
rect 111430 328170 111498 328226
rect 111554 328170 111622 328226
rect 111678 328170 115958 328226
rect 116014 328170 116082 328226
rect 116138 328170 146678 328226
rect 146734 328170 146802 328226
rect 146858 328170 177398 328226
rect 177454 328170 177522 328226
rect 177578 328170 208118 328226
rect 208174 328170 208242 328226
rect 208298 328170 238838 328226
rect 238894 328170 238962 328226
rect 239018 328170 269558 328226
rect 269614 328170 269682 328226
rect 269738 328170 300278 328226
rect 300334 328170 300402 328226
rect 300458 328170 330998 328226
rect 331054 328170 331122 328226
rect 331178 328170 361718 328226
rect 361774 328170 361842 328226
rect 361898 328170 392438 328226
rect 392494 328170 392562 328226
rect 392618 328170 423158 328226
rect 423214 328170 423282 328226
rect 423338 328170 453878 328226
rect 453934 328170 454002 328226
rect 454058 328170 484598 328226
rect 484654 328170 484722 328226
rect 484778 328170 515318 328226
rect 515374 328170 515442 328226
rect 515498 328170 546038 328226
rect 546094 328170 546162 328226
rect 546218 328170 561250 328226
rect 561306 328170 561374 328226
rect 561430 328170 561498 328226
rect 561554 328170 561622 328226
rect 561678 328170 579250 328226
rect 579306 328170 579374 328226
rect 579430 328170 579498 328226
rect 579554 328170 579622 328226
rect 579678 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597980 328226
rect -1916 328102 597980 328170
rect -1916 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 3250 328102
rect 3306 328046 3374 328102
rect 3430 328046 3498 328102
rect 3554 328046 3622 328102
rect 3678 328046 21250 328102
rect 21306 328046 21374 328102
rect 21430 328046 21498 328102
rect 21554 328046 21622 328102
rect 21678 328046 39250 328102
rect 39306 328046 39374 328102
rect 39430 328046 39498 328102
rect 39554 328046 39622 328102
rect 39678 328046 54518 328102
rect 54574 328046 54642 328102
rect 54698 328046 57250 328102
rect 57306 328046 57374 328102
rect 57430 328046 57498 328102
rect 57554 328046 57622 328102
rect 57678 328046 75250 328102
rect 75306 328046 75374 328102
rect 75430 328046 75498 328102
rect 75554 328046 75622 328102
rect 75678 328046 85238 328102
rect 85294 328046 85362 328102
rect 85418 328046 93250 328102
rect 93306 328046 93374 328102
rect 93430 328046 93498 328102
rect 93554 328046 93622 328102
rect 93678 328046 111250 328102
rect 111306 328046 111374 328102
rect 111430 328046 111498 328102
rect 111554 328046 111622 328102
rect 111678 328046 115958 328102
rect 116014 328046 116082 328102
rect 116138 328046 146678 328102
rect 146734 328046 146802 328102
rect 146858 328046 177398 328102
rect 177454 328046 177522 328102
rect 177578 328046 208118 328102
rect 208174 328046 208242 328102
rect 208298 328046 238838 328102
rect 238894 328046 238962 328102
rect 239018 328046 269558 328102
rect 269614 328046 269682 328102
rect 269738 328046 300278 328102
rect 300334 328046 300402 328102
rect 300458 328046 330998 328102
rect 331054 328046 331122 328102
rect 331178 328046 361718 328102
rect 361774 328046 361842 328102
rect 361898 328046 392438 328102
rect 392494 328046 392562 328102
rect 392618 328046 423158 328102
rect 423214 328046 423282 328102
rect 423338 328046 453878 328102
rect 453934 328046 454002 328102
rect 454058 328046 484598 328102
rect 484654 328046 484722 328102
rect 484778 328046 515318 328102
rect 515374 328046 515442 328102
rect 515498 328046 546038 328102
rect 546094 328046 546162 328102
rect 546218 328046 561250 328102
rect 561306 328046 561374 328102
rect 561430 328046 561498 328102
rect 561554 328046 561622 328102
rect 561678 328046 579250 328102
rect 579306 328046 579374 328102
rect 579430 328046 579498 328102
rect 579554 328046 579622 328102
rect 579678 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597980 328102
rect -1916 327978 597980 328046
rect -1916 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 3250 327978
rect 3306 327922 3374 327978
rect 3430 327922 3498 327978
rect 3554 327922 3622 327978
rect 3678 327922 21250 327978
rect 21306 327922 21374 327978
rect 21430 327922 21498 327978
rect 21554 327922 21622 327978
rect 21678 327922 39250 327978
rect 39306 327922 39374 327978
rect 39430 327922 39498 327978
rect 39554 327922 39622 327978
rect 39678 327922 54518 327978
rect 54574 327922 54642 327978
rect 54698 327922 57250 327978
rect 57306 327922 57374 327978
rect 57430 327922 57498 327978
rect 57554 327922 57622 327978
rect 57678 327922 75250 327978
rect 75306 327922 75374 327978
rect 75430 327922 75498 327978
rect 75554 327922 75622 327978
rect 75678 327922 85238 327978
rect 85294 327922 85362 327978
rect 85418 327922 93250 327978
rect 93306 327922 93374 327978
rect 93430 327922 93498 327978
rect 93554 327922 93622 327978
rect 93678 327922 111250 327978
rect 111306 327922 111374 327978
rect 111430 327922 111498 327978
rect 111554 327922 111622 327978
rect 111678 327922 115958 327978
rect 116014 327922 116082 327978
rect 116138 327922 146678 327978
rect 146734 327922 146802 327978
rect 146858 327922 177398 327978
rect 177454 327922 177522 327978
rect 177578 327922 208118 327978
rect 208174 327922 208242 327978
rect 208298 327922 238838 327978
rect 238894 327922 238962 327978
rect 239018 327922 269558 327978
rect 269614 327922 269682 327978
rect 269738 327922 300278 327978
rect 300334 327922 300402 327978
rect 300458 327922 330998 327978
rect 331054 327922 331122 327978
rect 331178 327922 361718 327978
rect 361774 327922 361842 327978
rect 361898 327922 392438 327978
rect 392494 327922 392562 327978
rect 392618 327922 423158 327978
rect 423214 327922 423282 327978
rect 423338 327922 453878 327978
rect 453934 327922 454002 327978
rect 454058 327922 484598 327978
rect 484654 327922 484722 327978
rect 484778 327922 515318 327978
rect 515374 327922 515442 327978
rect 515498 327922 546038 327978
rect 546094 327922 546162 327978
rect 546218 327922 561250 327978
rect 561306 327922 561374 327978
rect 561430 327922 561498 327978
rect 561554 327922 561622 327978
rect 561678 327922 579250 327978
rect 579306 327922 579374 327978
rect 579430 327922 579498 327978
rect 579554 327922 579622 327978
rect 579678 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597980 327978
rect -1916 327826 597980 327922
rect -1916 316350 597980 316446
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 6970 316350
rect 7026 316294 7094 316350
rect 7150 316294 7218 316350
rect 7274 316294 7342 316350
rect 7398 316294 24970 316350
rect 25026 316294 25094 316350
rect 25150 316294 25218 316350
rect 25274 316294 25342 316350
rect 25398 316294 42970 316350
rect 43026 316294 43094 316350
rect 43150 316294 43218 316350
rect 43274 316294 43342 316350
rect 43398 316294 60970 316350
rect 61026 316294 61094 316350
rect 61150 316294 61218 316350
rect 61274 316294 61342 316350
rect 61398 316294 69878 316350
rect 69934 316294 70002 316350
rect 70058 316294 78970 316350
rect 79026 316294 79094 316350
rect 79150 316294 79218 316350
rect 79274 316294 79342 316350
rect 79398 316294 96970 316350
rect 97026 316294 97094 316350
rect 97150 316294 97218 316350
rect 97274 316294 97342 316350
rect 97398 316294 100598 316350
rect 100654 316294 100722 316350
rect 100778 316294 131318 316350
rect 131374 316294 131442 316350
rect 131498 316294 162038 316350
rect 162094 316294 162162 316350
rect 162218 316294 192758 316350
rect 192814 316294 192882 316350
rect 192938 316294 223478 316350
rect 223534 316294 223602 316350
rect 223658 316294 254198 316350
rect 254254 316294 254322 316350
rect 254378 316294 284918 316350
rect 284974 316294 285042 316350
rect 285098 316294 315638 316350
rect 315694 316294 315762 316350
rect 315818 316294 346358 316350
rect 346414 316294 346482 316350
rect 346538 316294 377078 316350
rect 377134 316294 377202 316350
rect 377258 316294 407798 316350
rect 407854 316294 407922 316350
rect 407978 316294 438518 316350
rect 438574 316294 438642 316350
rect 438698 316294 469238 316350
rect 469294 316294 469362 316350
rect 469418 316294 499958 316350
rect 500014 316294 500082 316350
rect 500138 316294 530678 316350
rect 530734 316294 530802 316350
rect 530858 316294 564970 316350
rect 565026 316294 565094 316350
rect 565150 316294 565218 316350
rect 565274 316294 565342 316350
rect 565398 316294 582970 316350
rect 583026 316294 583094 316350
rect 583150 316294 583218 316350
rect 583274 316294 583342 316350
rect 583398 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect -1916 316226 597980 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 6970 316226
rect 7026 316170 7094 316226
rect 7150 316170 7218 316226
rect 7274 316170 7342 316226
rect 7398 316170 24970 316226
rect 25026 316170 25094 316226
rect 25150 316170 25218 316226
rect 25274 316170 25342 316226
rect 25398 316170 42970 316226
rect 43026 316170 43094 316226
rect 43150 316170 43218 316226
rect 43274 316170 43342 316226
rect 43398 316170 60970 316226
rect 61026 316170 61094 316226
rect 61150 316170 61218 316226
rect 61274 316170 61342 316226
rect 61398 316170 69878 316226
rect 69934 316170 70002 316226
rect 70058 316170 78970 316226
rect 79026 316170 79094 316226
rect 79150 316170 79218 316226
rect 79274 316170 79342 316226
rect 79398 316170 96970 316226
rect 97026 316170 97094 316226
rect 97150 316170 97218 316226
rect 97274 316170 97342 316226
rect 97398 316170 100598 316226
rect 100654 316170 100722 316226
rect 100778 316170 131318 316226
rect 131374 316170 131442 316226
rect 131498 316170 162038 316226
rect 162094 316170 162162 316226
rect 162218 316170 192758 316226
rect 192814 316170 192882 316226
rect 192938 316170 223478 316226
rect 223534 316170 223602 316226
rect 223658 316170 254198 316226
rect 254254 316170 254322 316226
rect 254378 316170 284918 316226
rect 284974 316170 285042 316226
rect 285098 316170 315638 316226
rect 315694 316170 315762 316226
rect 315818 316170 346358 316226
rect 346414 316170 346482 316226
rect 346538 316170 377078 316226
rect 377134 316170 377202 316226
rect 377258 316170 407798 316226
rect 407854 316170 407922 316226
rect 407978 316170 438518 316226
rect 438574 316170 438642 316226
rect 438698 316170 469238 316226
rect 469294 316170 469362 316226
rect 469418 316170 499958 316226
rect 500014 316170 500082 316226
rect 500138 316170 530678 316226
rect 530734 316170 530802 316226
rect 530858 316170 564970 316226
rect 565026 316170 565094 316226
rect 565150 316170 565218 316226
rect 565274 316170 565342 316226
rect 565398 316170 582970 316226
rect 583026 316170 583094 316226
rect 583150 316170 583218 316226
rect 583274 316170 583342 316226
rect 583398 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect -1916 316102 597980 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 6970 316102
rect 7026 316046 7094 316102
rect 7150 316046 7218 316102
rect 7274 316046 7342 316102
rect 7398 316046 24970 316102
rect 25026 316046 25094 316102
rect 25150 316046 25218 316102
rect 25274 316046 25342 316102
rect 25398 316046 42970 316102
rect 43026 316046 43094 316102
rect 43150 316046 43218 316102
rect 43274 316046 43342 316102
rect 43398 316046 60970 316102
rect 61026 316046 61094 316102
rect 61150 316046 61218 316102
rect 61274 316046 61342 316102
rect 61398 316046 69878 316102
rect 69934 316046 70002 316102
rect 70058 316046 78970 316102
rect 79026 316046 79094 316102
rect 79150 316046 79218 316102
rect 79274 316046 79342 316102
rect 79398 316046 96970 316102
rect 97026 316046 97094 316102
rect 97150 316046 97218 316102
rect 97274 316046 97342 316102
rect 97398 316046 100598 316102
rect 100654 316046 100722 316102
rect 100778 316046 131318 316102
rect 131374 316046 131442 316102
rect 131498 316046 162038 316102
rect 162094 316046 162162 316102
rect 162218 316046 192758 316102
rect 192814 316046 192882 316102
rect 192938 316046 223478 316102
rect 223534 316046 223602 316102
rect 223658 316046 254198 316102
rect 254254 316046 254322 316102
rect 254378 316046 284918 316102
rect 284974 316046 285042 316102
rect 285098 316046 315638 316102
rect 315694 316046 315762 316102
rect 315818 316046 346358 316102
rect 346414 316046 346482 316102
rect 346538 316046 377078 316102
rect 377134 316046 377202 316102
rect 377258 316046 407798 316102
rect 407854 316046 407922 316102
rect 407978 316046 438518 316102
rect 438574 316046 438642 316102
rect 438698 316046 469238 316102
rect 469294 316046 469362 316102
rect 469418 316046 499958 316102
rect 500014 316046 500082 316102
rect 500138 316046 530678 316102
rect 530734 316046 530802 316102
rect 530858 316046 564970 316102
rect 565026 316046 565094 316102
rect 565150 316046 565218 316102
rect 565274 316046 565342 316102
rect 565398 316046 582970 316102
rect 583026 316046 583094 316102
rect 583150 316046 583218 316102
rect 583274 316046 583342 316102
rect 583398 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect -1916 315978 597980 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 6970 315978
rect 7026 315922 7094 315978
rect 7150 315922 7218 315978
rect 7274 315922 7342 315978
rect 7398 315922 24970 315978
rect 25026 315922 25094 315978
rect 25150 315922 25218 315978
rect 25274 315922 25342 315978
rect 25398 315922 42970 315978
rect 43026 315922 43094 315978
rect 43150 315922 43218 315978
rect 43274 315922 43342 315978
rect 43398 315922 60970 315978
rect 61026 315922 61094 315978
rect 61150 315922 61218 315978
rect 61274 315922 61342 315978
rect 61398 315922 69878 315978
rect 69934 315922 70002 315978
rect 70058 315922 78970 315978
rect 79026 315922 79094 315978
rect 79150 315922 79218 315978
rect 79274 315922 79342 315978
rect 79398 315922 96970 315978
rect 97026 315922 97094 315978
rect 97150 315922 97218 315978
rect 97274 315922 97342 315978
rect 97398 315922 100598 315978
rect 100654 315922 100722 315978
rect 100778 315922 131318 315978
rect 131374 315922 131442 315978
rect 131498 315922 162038 315978
rect 162094 315922 162162 315978
rect 162218 315922 192758 315978
rect 192814 315922 192882 315978
rect 192938 315922 223478 315978
rect 223534 315922 223602 315978
rect 223658 315922 254198 315978
rect 254254 315922 254322 315978
rect 254378 315922 284918 315978
rect 284974 315922 285042 315978
rect 285098 315922 315638 315978
rect 315694 315922 315762 315978
rect 315818 315922 346358 315978
rect 346414 315922 346482 315978
rect 346538 315922 377078 315978
rect 377134 315922 377202 315978
rect 377258 315922 407798 315978
rect 407854 315922 407922 315978
rect 407978 315922 438518 315978
rect 438574 315922 438642 315978
rect 438698 315922 469238 315978
rect 469294 315922 469362 315978
rect 469418 315922 499958 315978
rect 500014 315922 500082 315978
rect 500138 315922 530678 315978
rect 530734 315922 530802 315978
rect 530858 315922 564970 315978
rect 565026 315922 565094 315978
rect 565150 315922 565218 315978
rect 565274 315922 565342 315978
rect 565398 315922 582970 315978
rect 583026 315922 583094 315978
rect 583150 315922 583218 315978
rect 583274 315922 583342 315978
rect 583398 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect -1916 315826 597980 315922
rect -1916 310350 597980 310446
rect -1916 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 3250 310350
rect 3306 310294 3374 310350
rect 3430 310294 3498 310350
rect 3554 310294 3622 310350
rect 3678 310294 21250 310350
rect 21306 310294 21374 310350
rect 21430 310294 21498 310350
rect 21554 310294 21622 310350
rect 21678 310294 39250 310350
rect 39306 310294 39374 310350
rect 39430 310294 39498 310350
rect 39554 310294 39622 310350
rect 39678 310294 54518 310350
rect 54574 310294 54642 310350
rect 54698 310294 57250 310350
rect 57306 310294 57374 310350
rect 57430 310294 57498 310350
rect 57554 310294 57622 310350
rect 57678 310294 75250 310350
rect 75306 310294 75374 310350
rect 75430 310294 75498 310350
rect 75554 310294 75622 310350
rect 75678 310294 85238 310350
rect 85294 310294 85362 310350
rect 85418 310294 93250 310350
rect 93306 310294 93374 310350
rect 93430 310294 93498 310350
rect 93554 310294 93622 310350
rect 93678 310294 111250 310350
rect 111306 310294 111374 310350
rect 111430 310294 111498 310350
rect 111554 310294 111622 310350
rect 111678 310294 115958 310350
rect 116014 310294 116082 310350
rect 116138 310294 146678 310350
rect 146734 310294 146802 310350
rect 146858 310294 177398 310350
rect 177454 310294 177522 310350
rect 177578 310294 208118 310350
rect 208174 310294 208242 310350
rect 208298 310294 238838 310350
rect 238894 310294 238962 310350
rect 239018 310294 269558 310350
rect 269614 310294 269682 310350
rect 269738 310294 300278 310350
rect 300334 310294 300402 310350
rect 300458 310294 330998 310350
rect 331054 310294 331122 310350
rect 331178 310294 361718 310350
rect 361774 310294 361842 310350
rect 361898 310294 392438 310350
rect 392494 310294 392562 310350
rect 392618 310294 423158 310350
rect 423214 310294 423282 310350
rect 423338 310294 453878 310350
rect 453934 310294 454002 310350
rect 454058 310294 484598 310350
rect 484654 310294 484722 310350
rect 484778 310294 515318 310350
rect 515374 310294 515442 310350
rect 515498 310294 546038 310350
rect 546094 310294 546162 310350
rect 546218 310294 561250 310350
rect 561306 310294 561374 310350
rect 561430 310294 561498 310350
rect 561554 310294 561622 310350
rect 561678 310294 579250 310350
rect 579306 310294 579374 310350
rect 579430 310294 579498 310350
rect 579554 310294 579622 310350
rect 579678 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597980 310350
rect -1916 310226 597980 310294
rect -1916 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 3250 310226
rect 3306 310170 3374 310226
rect 3430 310170 3498 310226
rect 3554 310170 3622 310226
rect 3678 310170 21250 310226
rect 21306 310170 21374 310226
rect 21430 310170 21498 310226
rect 21554 310170 21622 310226
rect 21678 310170 39250 310226
rect 39306 310170 39374 310226
rect 39430 310170 39498 310226
rect 39554 310170 39622 310226
rect 39678 310170 54518 310226
rect 54574 310170 54642 310226
rect 54698 310170 57250 310226
rect 57306 310170 57374 310226
rect 57430 310170 57498 310226
rect 57554 310170 57622 310226
rect 57678 310170 75250 310226
rect 75306 310170 75374 310226
rect 75430 310170 75498 310226
rect 75554 310170 75622 310226
rect 75678 310170 85238 310226
rect 85294 310170 85362 310226
rect 85418 310170 93250 310226
rect 93306 310170 93374 310226
rect 93430 310170 93498 310226
rect 93554 310170 93622 310226
rect 93678 310170 111250 310226
rect 111306 310170 111374 310226
rect 111430 310170 111498 310226
rect 111554 310170 111622 310226
rect 111678 310170 115958 310226
rect 116014 310170 116082 310226
rect 116138 310170 146678 310226
rect 146734 310170 146802 310226
rect 146858 310170 177398 310226
rect 177454 310170 177522 310226
rect 177578 310170 208118 310226
rect 208174 310170 208242 310226
rect 208298 310170 238838 310226
rect 238894 310170 238962 310226
rect 239018 310170 269558 310226
rect 269614 310170 269682 310226
rect 269738 310170 300278 310226
rect 300334 310170 300402 310226
rect 300458 310170 330998 310226
rect 331054 310170 331122 310226
rect 331178 310170 361718 310226
rect 361774 310170 361842 310226
rect 361898 310170 392438 310226
rect 392494 310170 392562 310226
rect 392618 310170 423158 310226
rect 423214 310170 423282 310226
rect 423338 310170 453878 310226
rect 453934 310170 454002 310226
rect 454058 310170 484598 310226
rect 484654 310170 484722 310226
rect 484778 310170 515318 310226
rect 515374 310170 515442 310226
rect 515498 310170 546038 310226
rect 546094 310170 546162 310226
rect 546218 310170 561250 310226
rect 561306 310170 561374 310226
rect 561430 310170 561498 310226
rect 561554 310170 561622 310226
rect 561678 310170 579250 310226
rect 579306 310170 579374 310226
rect 579430 310170 579498 310226
rect 579554 310170 579622 310226
rect 579678 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597980 310226
rect -1916 310102 597980 310170
rect -1916 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 3250 310102
rect 3306 310046 3374 310102
rect 3430 310046 3498 310102
rect 3554 310046 3622 310102
rect 3678 310046 21250 310102
rect 21306 310046 21374 310102
rect 21430 310046 21498 310102
rect 21554 310046 21622 310102
rect 21678 310046 39250 310102
rect 39306 310046 39374 310102
rect 39430 310046 39498 310102
rect 39554 310046 39622 310102
rect 39678 310046 54518 310102
rect 54574 310046 54642 310102
rect 54698 310046 57250 310102
rect 57306 310046 57374 310102
rect 57430 310046 57498 310102
rect 57554 310046 57622 310102
rect 57678 310046 75250 310102
rect 75306 310046 75374 310102
rect 75430 310046 75498 310102
rect 75554 310046 75622 310102
rect 75678 310046 85238 310102
rect 85294 310046 85362 310102
rect 85418 310046 93250 310102
rect 93306 310046 93374 310102
rect 93430 310046 93498 310102
rect 93554 310046 93622 310102
rect 93678 310046 111250 310102
rect 111306 310046 111374 310102
rect 111430 310046 111498 310102
rect 111554 310046 111622 310102
rect 111678 310046 115958 310102
rect 116014 310046 116082 310102
rect 116138 310046 146678 310102
rect 146734 310046 146802 310102
rect 146858 310046 177398 310102
rect 177454 310046 177522 310102
rect 177578 310046 208118 310102
rect 208174 310046 208242 310102
rect 208298 310046 238838 310102
rect 238894 310046 238962 310102
rect 239018 310046 269558 310102
rect 269614 310046 269682 310102
rect 269738 310046 300278 310102
rect 300334 310046 300402 310102
rect 300458 310046 330998 310102
rect 331054 310046 331122 310102
rect 331178 310046 361718 310102
rect 361774 310046 361842 310102
rect 361898 310046 392438 310102
rect 392494 310046 392562 310102
rect 392618 310046 423158 310102
rect 423214 310046 423282 310102
rect 423338 310046 453878 310102
rect 453934 310046 454002 310102
rect 454058 310046 484598 310102
rect 484654 310046 484722 310102
rect 484778 310046 515318 310102
rect 515374 310046 515442 310102
rect 515498 310046 546038 310102
rect 546094 310046 546162 310102
rect 546218 310046 561250 310102
rect 561306 310046 561374 310102
rect 561430 310046 561498 310102
rect 561554 310046 561622 310102
rect 561678 310046 579250 310102
rect 579306 310046 579374 310102
rect 579430 310046 579498 310102
rect 579554 310046 579622 310102
rect 579678 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597980 310102
rect -1916 309978 597980 310046
rect -1916 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 3250 309978
rect 3306 309922 3374 309978
rect 3430 309922 3498 309978
rect 3554 309922 3622 309978
rect 3678 309922 21250 309978
rect 21306 309922 21374 309978
rect 21430 309922 21498 309978
rect 21554 309922 21622 309978
rect 21678 309922 39250 309978
rect 39306 309922 39374 309978
rect 39430 309922 39498 309978
rect 39554 309922 39622 309978
rect 39678 309922 54518 309978
rect 54574 309922 54642 309978
rect 54698 309922 57250 309978
rect 57306 309922 57374 309978
rect 57430 309922 57498 309978
rect 57554 309922 57622 309978
rect 57678 309922 75250 309978
rect 75306 309922 75374 309978
rect 75430 309922 75498 309978
rect 75554 309922 75622 309978
rect 75678 309922 85238 309978
rect 85294 309922 85362 309978
rect 85418 309922 93250 309978
rect 93306 309922 93374 309978
rect 93430 309922 93498 309978
rect 93554 309922 93622 309978
rect 93678 309922 111250 309978
rect 111306 309922 111374 309978
rect 111430 309922 111498 309978
rect 111554 309922 111622 309978
rect 111678 309922 115958 309978
rect 116014 309922 116082 309978
rect 116138 309922 146678 309978
rect 146734 309922 146802 309978
rect 146858 309922 177398 309978
rect 177454 309922 177522 309978
rect 177578 309922 208118 309978
rect 208174 309922 208242 309978
rect 208298 309922 238838 309978
rect 238894 309922 238962 309978
rect 239018 309922 269558 309978
rect 269614 309922 269682 309978
rect 269738 309922 300278 309978
rect 300334 309922 300402 309978
rect 300458 309922 330998 309978
rect 331054 309922 331122 309978
rect 331178 309922 361718 309978
rect 361774 309922 361842 309978
rect 361898 309922 392438 309978
rect 392494 309922 392562 309978
rect 392618 309922 423158 309978
rect 423214 309922 423282 309978
rect 423338 309922 453878 309978
rect 453934 309922 454002 309978
rect 454058 309922 484598 309978
rect 484654 309922 484722 309978
rect 484778 309922 515318 309978
rect 515374 309922 515442 309978
rect 515498 309922 546038 309978
rect 546094 309922 546162 309978
rect 546218 309922 561250 309978
rect 561306 309922 561374 309978
rect 561430 309922 561498 309978
rect 561554 309922 561622 309978
rect 561678 309922 579250 309978
rect 579306 309922 579374 309978
rect 579430 309922 579498 309978
rect 579554 309922 579622 309978
rect 579678 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597980 309978
rect -1916 309826 597980 309922
rect -1916 298350 597980 298446
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 6970 298350
rect 7026 298294 7094 298350
rect 7150 298294 7218 298350
rect 7274 298294 7342 298350
rect 7398 298294 24970 298350
rect 25026 298294 25094 298350
rect 25150 298294 25218 298350
rect 25274 298294 25342 298350
rect 25398 298294 42970 298350
rect 43026 298294 43094 298350
rect 43150 298294 43218 298350
rect 43274 298294 43342 298350
rect 43398 298294 60970 298350
rect 61026 298294 61094 298350
rect 61150 298294 61218 298350
rect 61274 298294 61342 298350
rect 61398 298294 69878 298350
rect 69934 298294 70002 298350
rect 70058 298294 78970 298350
rect 79026 298294 79094 298350
rect 79150 298294 79218 298350
rect 79274 298294 79342 298350
rect 79398 298294 96970 298350
rect 97026 298294 97094 298350
rect 97150 298294 97218 298350
rect 97274 298294 97342 298350
rect 97398 298294 100598 298350
rect 100654 298294 100722 298350
rect 100778 298294 131318 298350
rect 131374 298294 131442 298350
rect 131498 298294 162038 298350
rect 162094 298294 162162 298350
rect 162218 298294 192758 298350
rect 192814 298294 192882 298350
rect 192938 298294 223478 298350
rect 223534 298294 223602 298350
rect 223658 298294 254198 298350
rect 254254 298294 254322 298350
rect 254378 298294 284918 298350
rect 284974 298294 285042 298350
rect 285098 298294 315638 298350
rect 315694 298294 315762 298350
rect 315818 298294 346358 298350
rect 346414 298294 346482 298350
rect 346538 298294 377078 298350
rect 377134 298294 377202 298350
rect 377258 298294 407798 298350
rect 407854 298294 407922 298350
rect 407978 298294 438518 298350
rect 438574 298294 438642 298350
rect 438698 298294 469238 298350
rect 469294 298294 469362 298350
rect 469418 298294 499958 298350
rect 500014 298294 500082 298350
rect 500138 298294 530678 298350
rect 530734 298294 530802 298350
rect 530858 298294 564970 298350
rect 565026 298294 565094 298350
rect 565150 298294 565218 298350
rect 565274 298294 565342 298350
rect 565398 298294 582970 298350
rect 583026 298294 583094 298350
rect 583150 298294 583218 298350
rect 583274 298294 583342 298350
rect 583398 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect -1916 298226 597980 298294
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 6970 298226
rect 7026 298170 7094 298226
rect 7150 298170 7218 298226
rect 7274 298170 7342 298226
rect 7398 298170 24970 298226
rect 25026 298170 25094 298226
rect 25150 298170 25218 298226
rect 25274 298170 25342 298226
rect 25398 298170 42970 298226
rect 43026 298170 43094 298226
rect 43150 298170 43218 298226
rect 43274 298170 43342 298226
rect 43398 298170 60970 298226
rect 61026 298170 61094 298226
rect 61150 298170 61218 298226
rect 61274 298170 61342 298226
rect 61398 298170 69878 298226
rect 69934 298170 70002 298226
rect 70058 298170 78970 298226
rect 79026 298170 79094 298226
rect 79150 298170 79218 298226
rect 79274 298170 79342 298226
rect 79398 298170 96970 298226
rect 97026 298170 97094 298226
rect 97150 298170 97218 298226
rect 97274 298170 97342 298226
rect 97398 298170 100598 298226
rect 100654 298170 100722 298226
rect 100778 298170 131318 298226
rect 131374 298170 131442 298226
rect 131498 298170 162038 298226
rect 162094 298170 162162 298226
rect 162218 298170 192758 298226
rect 192814 298170 192882 298226
rect 192938 298170 223478 298226
rect 223534 298170 223602 298226
rect 223658 298170 254198 298226
rect 254254 298170 254322 298226
rect 254378 298170 284918 298226
rect 284974 298170 285042 298226
rect 285098 298170 315638 298226
rect 315694 298170 315762 298226
rect 315818 298170 346358 298226
rect 346414 298170 346482 298226
rect 346538 298170 377078 298226
rect 377134 298170 377202 298226
rect 377258 298170 407798 298226
rect 407854 298170 407922 298226
rect 407978 298170 438518 298226
rect 438574 298170 438642 298226
rect 438698 298170 469238 298226
rect 469294 298170 469362 298226
rect 469418 298170 499958 298226
rect 500014 298170 500082 298226
rect 500138 298170 530678 298226
rect 530734 298170 530802 298226
rect 530858 298170 564970 298226
rect 565026 298170 565094 298226
rect 565150 298170 565218 298226
rect 565274 298170 565342 298226
rect 565398 298170 582970 298226
rect 583026 298170 583094 298226
rect 583150 298170 583218 298226
rect 583274 298170 583342 298226
rect 583398 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect -1916 298102 597980 298170
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 6970 298102
rect 7026 298046 7094 298102
rect 7150 298046 7218 298102
rect 7274 298046 7342 298102
rect 7398 298046 24970 298102
rect 25026 298046 25094 298102
rect 25150 298046 25218 298102
rect 25274 298046 25342 298102
rect 25398 298046 42970 298102
rect 43026 298046 43094 298102
rect 43150 298046 43218 298102
rect 43274 298046 43342 298102
rect 43398 298046 60970 298102
rect 61026 298046 61094 298102
rect 61150 298046 61218 298102
rect 61274 298046 61342 298102
rect 61398 298046 69878 298102
rect 69934 298046 70002 298102
rect 70058 298046 78970 298102
rect 79026 298046 79094 298102
rect 79150 298046 79218 298102
rect 79274 298046 79342 298102
rect 79398 298046 96970 298102
rect 97026 298046 97094 298102
rect 97150 298046 97218 298102
rect 97274 298046 97342 298102
rect 97398 298046 100598 298102
rect 100654 298046 100722 298102
rect 100778 298046 131318 298102
rect 131374 298046 131442 298102
rect 131498 298046 162038 298102
rect 162094 298046 162162 298102
rect 162218 298046 192758 298102
rect 192814 298046 192882 298102
rect 192938 298046 223478 298102
rect 223534 298046 223602 298102
rect 223658 298046 254198 298102
rect 254254 298046 254322 298102
rect 254378 298046 284918 298102
rect 284974 298046 285042 298102
rect 285098 298046 315638 298102
rect 315694 298046 315762 298102
rect 315818 298046 346358 298102
rect 346414 298046 346482 298102
rect 346538 298046 377078 298102
rect 377134 298046 377202 298102
rect 377258 298046 407798 298102
rect 407854 298046 407922 298102
rect 407978 298046 438518 298102
rect 438574 298046 438642 298102
rect 438698 298046 469238 298102
rect 469294 298046 469362 298102
rect 469418 298046 499958 298102
rect 500014 298046 500082 298102
rect 500138 298046 530678 298102
rect 530734 298046 530802 298102
rect 530858 298046 564970 298102
rect 565026 298046 565094 298102
rect 565150 298046 565218 298102
rect 565274 298046 565342 298102
rect 565398 298046 582970 298102
rect 583026 298046 583094 298102
rect 583150 298046 583218 298102
rect 583274 298046 583342 298102
rect 583398 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect -1916 297978 597980 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 6970 297978
rect 7026 297922 7094 297978
rect 7150 297922 7218 297978
rect 7274 297922 7342 297978
rect 7398 297922 24970 297978
rect 25026 297922 25094 297978
rect 25150 297922 25218 297978
rect 25274 297922 25342 297978
rect 25398 297922 42970 297978
rect 43026 297922 43094 297978
rect 43150 297922 43218 297978
rect 43274 297922 43342 297978
rect 43398 297922 60970 297978
rect 61026 297922 61094 297978
rect 61150 297922 61218 297978
rect 61274 297922 61342 297978
rect 61398 297922 69878 297978
rect 69934 297922 70002 297978
rect 70058 297922 78970 297978
rect 79026 297922 79094 297978
rect 79150 297922 79218 297978
rect 79274 297922 79342 297978
rect 79398 297922 96970 297978
rect 97026 297922 97094 297978
rect 97150 297922 97218 297978
rect 97274 297922 97342 297978
rect 97398 297922 100598 297978
rect 100654 297922 100722 297978
rect 100778 297922 131318 297978
rect 131374 297922 131442 297978
rect 131498 297922 162038 297978
rect 162094 297922 162162 297978
rect 162218 297922 192758 297978
rect 192814 297922 192882 297978
rect 192938 297922 223478 297978
rect 223534 297922 223602 297978
rect 223658 297922 254198 297978
rect 254254 297922 254322 297978
rect 254378 297922 284918 297978
rect 284974 297922 285042 297978
rect 285098 297922 315638 297978
rect 315694 297922 315762 297978
rect 315818 297922 346358 297978
rect 346414 297922 346482 297978
rect 346538 297922 377078 297978
rect 377134 297922 377202 297978
rect 377258 297922 407798 297978
rect 407854 297922 407922 297978
rect 407978 297922 438518 297978
rect 438574 297922 438642 297978
rect 438698 297922 469238 297978
rect 469294 297922 469362 297978
rect 469418 297922 499958 297978
rect 500014 297922 500082 297978
rect 500138 297922 530678 297978
rect 530734 297922 530802 297978
rect 530858 297922 564970 297978
rect 565026 297922 565094 297978
rect 565150 297922 565218 297978
rect 565274 297922 565342 297978
rect 565398 297922 582970 297978
rect 583026 297922 583094 297978
rect 583150 297922 583218 297978
rect 583274 297922 583342 297978
rect 583398 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect -1916 297826 597980 297922
rect -1916 292350 597980 292446
rect -1916 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 3250 292350
rect 3306 292294 3374 292350
rect 3430 292294 3498 292350
rect 3554 292294 3622 292350
rect 3678 292294 21250 292350
rect 21306 292294 21374 292350
rect 21430 292294 21498 292350
rect 21554 292294 21622 292350
rect 21678 292294 39250 292350
rect 39306 292294 39374 292350
rect 39430 292294 39498 292350
rect 39554 292294 39622 292350
rect 39678 292294 54518 292350
rect 54574 292294 54642 292350
rect 54698 292294 57250 292350
rect 57306 292294 57374 292350
rect 57430 292294 57498 292350
rect 57554 292294 57622 292350
rect 57678 292294 75250 292350
rect 75306 292294 75374 292350
rect 75430 292294 75498 292350
rect 75554 292294 75622 292350
rect 75678 292294 85238 292350
rect 85294 292294 85362 292350
rect 85418 292294 93250 292350
rect 93306 292294 93374 292350
rect 93430 292294 93498 292350
rect 93554 292294 93622 292350
rect 93678 292294 111250 292350
rect 111306 292294 111374 292350
rect 111430 292294 111498 292350
rect 111554 292294 111622 292350
rect 111678 292294 115958 292350
rect 116014 292294 116082 292350
rect 116138 292294 146678 292350
rect 146734 292294 146802 292350
rect 146858 292294 177398 292350
rect 177454 292294 177522 292350
rect 177578 292294 208118 292350
rect 208174 292294 208242 292350
rect 208298 292294 238838 292350
rect 238894 292294 238962 292350
rect 239018 292294 269558 292350
rect 269614 292294 269682 292350
rect 269738 292294 300278 292350
rect 300334 292294 300402 292350
rect 300458 292294 330998 292350
rect 331054 292294 331122 292350
rect 331178 292294 361718 292350
rect 361774 292294 361842 292350
rect 361898 292294 392438 292350
rect 392494 292294 392562 292350
rect 392618 292294 423158 292350
rect 423214 292294 423282 292350
rect 423338 292294 453878 292350
rect 453934 292294 454002 292350
rect 454058 292294 484598 292350
rect 484654 292294 484722 292350
rect 484778 292294 515318 292350
rect 515374 292294 515442 292350
rect 515498 292294 546038 292350
rect 546094 292294 546162 292350
rect 546218 292294 561250 292350
rect 561306 292294 561374 292350
rect 561430 292294 561498 292350
rect 561554 292294 561622 292350
rect 561678 292294 579250 292350
rect 579306 292294 579374 292350
rect 579430 292294 579498 292350
rect 579554 292294 579622 292350
rect 579678 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597980 292350
rect -1916 292226 597980 292294
rect -1916 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 3250 292226
rect 3306 292170 3374 292226
rect 3430 292170 3498 292226
rect 3554 292170 3622 292226
rect 3678 292170 21250 292226
rect 21306 292170 21374 292226
rect 21430 292170 21498 292226
rect 21554 292170 21622 292226
rect 21678 292170 39250 292226
rect 39306 292170 39374 292226
rect 39430 292170 39498 292226
rect 39554 292170 39622 292226
rect 39678 292170 54518 292226
rect 54574 292170 54642 292226
rect 54698 292170 57250 292226
rect 57306 292170 57374 292226
rect 57430 292170 57498 292226
rect 57554 292170 57622 292226
rect 57678 292170 75250 292226
rect 75306 292170 75374 292226
rect 75430 292170 75498 292226
rect 75554 292170 75622 292226
rect 75678 292170 85238 292226
rect 85294 292170 85362 292226
rect 85418 292170 93250 292226
rect 93306 292170 93374 292226
rect 93430 292170 93498 292226
rect 93554 292170 93622 292226
rect 93678 292170 111250 292226
rect 111306 292170 111374 292226
rect 111430 292170 111498 292226
rect 111554 292170 111622 292226
rect 111678 292170 115958 292226
rect 116014 292170 116082 292226
rect 116138 292170 146678 292226
rect 146734 292170 146802 292226
rect 146858 292170 177398 292226
rect 177454 292170 177522 292226
rect 177578 292170 208118 292226
rect 208174 292170 208242 292226
rect 208298 292170 238838 292226
rect 238894 292170 238962 292226
rect 239018 292170 269558 292226
rect 269614 292170 269682 292226
rect 269738 292170 300278 292226
rect 300334 292170 300402 292226
rect 300458 292170 330998 292226
rect 331054 292170 331122 292226
rect 331178 292170 361718 292226
rect 361774 292170 361842 292226
rect 361898 292170 392438 292226
rect 392494 292170 392562 292226
rect 392618 292170 423158 292226
rect 423214 292170 423282 292226
rect 423338 292170 453878 292226
rect 453934 292170 454002 292226
rect 454058 292170 484598 292226
rect 484654 292170 484722 292226
rect 484778 292170 515318 292226
rect 515374 292170 515442 292226
rect 515498 292170 546038 292226
rect 546094 292170 546162 292226
rect 546218 292170 561250 292226
rect 561306 292170 561374 292226
rect 561430 292170 561498 292226
rect 561554 292170 561622 292226
rect 561678 292170 579250 292226
rect 579306 292170 579374 292226
rect 579430 292170 579498 292226
rect 579554 292170 579622 292226
rect 579678 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597980 292226
rect -1916 292102 597980 292170
rect -1916 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 3250 292102
rect 3306 292046 3374 292102
rect 3430 292046 3498 292102
rect 3554 292046 3622 292102
rect 3678 292046 21250 292102
rect 21306 292046 21374 292102
rect 21430 292046 21498 292102
rect 21554 292046 21622 292102
rect 21678 292046 39250 292102
rect 39306 292046 39374 292102
rect 39430 292046 39498 292102
rect 39554 292046 39622 292102
rect 39678 292046 54518 292102
rect 54574 292046 54642 292102
rect 54698 292046 57250 292102
rect 57306 292046 57374 292102
rect 57430 292046 57498 292102
rect 57554 292046 57622 292102
rect 57678 292046 75250 292102
rect 75306 292046 75374 292102
rect 75430 292046 75498 292102
rect 75554 292046 75622 292102
rect 75678 292046 85238 292102
rect 85294 292046 85362 292102
rect 85418 292046 93250 292102
rect 93306 292046 93374 292102
rect 93430 292046 93498 292102
rect 93554 292046 93622 292102
rect 93678 292046 111250 292102
rect 111306 292046 111374 292102
rect 111430 292046 111498 292102
rect 111554 292046 111622 292102
rect 111678 292046 115958 292102
rect 116014 292046 116082 292102
rect 116138 292046 146678 292102
rect 146734 292046 146802 292102
rect 146858 292046 177398 292102
rect 177454 292046 177522 292102
rect 177578 292046 208118 292102
rect 208174 292046 208242 292102
rect 208298 292046 238838 292102
rect 238894 292046 238962 292102
rect 239018 292046 269558 292102
rect 269614 292046 269682 292102
rect 269738 292046 300278 292102
rect 300334 292046 300402 292102
rect 300458 292046 330998 292102
rect 331054 292046 331122 292102
rect 331178 292046 361718 292102
rect 361774 292046 361842 292102
rect 361898 292046 392438 292102
rect 392494 292046 392562 292102
rect 392618 292046 423158 292102
rect 423214 292046 423282 292102
rect 423338 292046 453878 292102
rect 453934 292046 454002 292102
rect 454058 292046 484598 292102
rect 484654 292046 484722 292102
rect 484778 292046 515318 292102
rect 515374 292046 515442 292102
rect 515498 292046 546038 292102
rect 546094 292046 546162 292102
rect 546218 292046 561250 292102
rect 561306 292046 561374 292102
rect 561430 292046 561498 292102
rect 561554 292046 561622 292102
rect 561678 292046 579250 292102
rect 579306 292046 579374 292102
rect 579430 292046 579498 292102
rect 579554 292046 579622 292102
rect 579678 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597980 292102
rect -1916 291978 597980 292046
rect -1916 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 3250 291978
rect 3306 291922 3374 291978
rect 3430 291922 3498 291978
rect 3554 291922 3622 291978
rect 3678 291922 21250 291978
rect 21306 291922 21374 291978
rect 21430 291922 21498 291978
rect 21554 291922 21622 291978
rect 21678 291922 39250 291978
rect 39306 291922 39374 291978
rect 39430 291922 39498 291978
rect 39554 291922 39622 291978
rect 39678 291922 54518 291978
rect 54574 291922 54642 291978
rect 54698 291922 57250 291978
rect 57306 291922 57374 291978
rect 57430 291922 57498 291978
rect 57554 291922 57622 291978
rect 57678 291922 75250 291978
rect 75306 291922 75374 291978
rect 75430 291922 75498 291978
rect 75554 291922 75622 291978
rect 75678 291922 85238 291978
rect 85294 291922 85362 291978
rect 85418 291922 93250 291978
rect 93306 291922 93374 291978
rect 93430 291922 93498 291978
rect 93554 291922 93622 291978
rect 93678 291922 111250 291978
rect 111306 291922 111374 291978
rect 111430 291922 111498 291978
rect 111554 291922 111622 291978
rect 111678 291922 115958 291978
rect 116014 291922 116082 291978
rect 116138 291922 146678 291978
rect 146734 291922 146802 291978
rect 146858 291922 177398 291978
rect 177454 291922 177522 291978
rect 177578 291922 208118 291978
rect 208174 291922 208242 291978
rect 208298 291922 238838 291978
rect 238894 291922 238962 291978
rect 239018 291922 269558 291978
rect 269614 291922 269682 291978
rect 269738 291922 300278 291978
rect 300334 291922 300402 291978
rect 300458 291922 330998 291978
rect 331054 291922 331122 291978
rect 331178 291922 361718 291978
rect 361774 291922 361842 291978
rect 361898 291922 392438 291978
rect 392494 291922 392562 291978
rect 392618 291922 423158 291978
rect 423214 291922 423282 291978
rect 423338 291922 453878 291978
rect 453934 291922 454002 291978
rect 454058 291922 484598 291978
rect 484654 291922 484722 291978
rect 484778 291922 515318 291978
rect 515374 291922 515442 291978
rect 515498 291922 546038 291978
rect 546094 291922 546162 291978
rect 546218 291922 561250 291978
rect 561306 291922 561374 291978
rect 561430 291922 561498 291978
rect 561554 291922 561622 291978
rect 561678 291922 579250 291978
rect 579306 291922 579374 291978
rect 579430 291922 579498 291978
rect 579554 291922 579622 291978
rect 579678 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597980 291978
rect -1916 291826 597980 291922
rect -1916 280350 597980 280446
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 6970 280350
rect 7026 280294 7094 280350
rect 7150 280294 7218 280350
rect 7274 280294 7342 280350
rect 7398 280294 24970 280350
rect 25026 280294 25094 280350
rect 25150 280294 25218 280350
rect 25274 280294 25342 280350
rect 25398 280294 42970 280350
rect 43026 280294 43094 280350
rect 43150 280294 43218 280350
rect 43274 280294 43342 280350
rect 43398 280294 60970 280350
rect 61026 280294 61094 280350
rect 61150 280294 61218 280350
rect 61274 280294 61342 280350
rect 61398 280294 69878 280350
rect 69934 280294 70002 280350
rect 70058 280294 78970 280350
rect 79026 280294 79094 280350
rect 79150 280294 79218 280350
rect 79274 280294 79342 280350
rect 79398 280294 96970 280350
rect 97026 280294 97094 280350
rect 97150 280294 97218 280350
rect 97274 280294 97342 280350
rect 97398 280294 100598 280350
rect 100654 280294 100722 280350
rect 100778 280294 131318 280350
rect 131374 280294 131442 280350
rect 131498 280294 162038 280350
rect 162094 280294 162162 280350
rect 162218 280294 192758 280350
rect 192814 280294 192882 280350
rect 192938 280294 223478 280350
rect 223534 280294 223602 280350
rect 223658 280294 254198 280350
rect 254254 280294 254322 280350
rect 254378 280294 284918 280350
rect 284974 280294 285042 280350
rect 285098 280294 315638 280350
rect 315694 280294 315762 280350
rect 315818 280294 346358 280350
rect 346414 280294 346482 280350
rect 346538 280294 377078 280350
rect 377134 280294 377202 280350
rect 377258 280294 407798 280350
rect 407854 280294 407922 280350
rect 407978 280294 438518 280350
rect 438574 280294 438642 280350
rect 438698 280294 469238 280350
rect 469294 280294 469362 280350
rect 469418 280294 499958 280350
rect 500014 280294 500082 280350
rect 500138 280294 530678 280350
rect 530734 280294 530802 280350
rect 530858 280294 564970 280350
rect 565026 280294 565094 280350
rect 565150 280294 565218 280350
rect 565274 280294 565342 280350
rect 565398 280294 582970 280350
rect 583026 280294 583094 280350
rect 583150 280294 583218 280350
rect 583274 280294 583342 280350
rect 583398 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect -1916 280226 597980 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 6970 280226
rect 7026 280170 7094 280226
rect 7150 280170 7218 280226
rect 7274 280170 7342 280226
rect 7398 280170 24970 280226
rect 25026 280170 25094 280226
rect 25150 280170 25218 280226
rect 25274 280170 25342 280226
rect 25398 280170 42970 280226
rect 43026 280170 43094 280226
rect 43150 280170 43218 280226
rect 43274 280170 43342 280226
rect 43398 280170 60970 280226
rect 61026 280170 61094 280226
rect 61150 280170 61218 280226
rect 61274 280170 61342 280226
rect 61398 280170 69878 280226
rect 69934 280170 70002 280226
rect 70058 280170 78970 280226
rect 79026 280170 79094 280226
rect 79150 280170 79218 280226
rect 79274 280170 79342 280226
rect 79398 280170 96970 280226
rect 97026 280170 97094 280226
rect 97150 280170 97218 280226
rect 97274 280170 97342 280226
rect 97398 280170 100598 280226
rect 100654 280170 100722 280226
rect 100778 280170 131318 280226
rect 131374 280170 131442 280226
rect 131498 280170 162038 280226
rect 162094 280170 162162 280226
rect 162218 280170 192758 280226
rect 192814 280170 192882 280226
rect 192938 280170 223478 280226
rect 223534 280170 223602 280226
rect 223658 280170 254198 280226
rect 254254 280170 254322 280226
rect 254378 280170 284918 280226
rect 284974 280170 285042 280226
rect 285098 280170 315638 280226
rect 315694 280170 315762 280226
rect 315818 280170 346358 280226
rect 346414 280170 346482 280226
rect 346538 280170 377078 280226
rect 377134 280170 377202 280226
rect 377258 280170 407798 280226
rect 407854 280170 407922 280226
rect 407978 280170 438518 280226
rect 438574 280170 438642 280226
rect 438698 280170 469238 280226
rect 469294 280170 469362 280226
rect 469418 280170 499958 280226
rect 500014 280170 500082 280226
rect 500138 280170 530678 280226
rect 530734 280170 530802 280226
rect 530858 280170 564970 280226
rect 565026 280170 565094 280226
rect 565150 280170 565218 280226
rect 565274 280170 565342 280226
rect 565398 280170 582970 280226
rect 583026 280170 583094 280226
rect 583150 280170 583218 280226
rect 583274 280170 583342 280226
rect 583398 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect -1916 280102 597980 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 6970 280102
rect 7026 280046 7094 280102
rect 7150 280046 7218 280102
rect 7274 280046 7342 280102
rect 7398 280046 24970 280102
rect 25026 280046 25094 280102
rect 25150 280046 25218 280102
rect 25274 280046 25342 280102
rect 25398 280046 42970 280102
rect 43026 280046 43094 280102
rect 43150 280046 43218 280102
rect 43274 280046 43342 280102
rect 43398 280046 60970 280102
rect 61026 280046 61094 280102
rect 61150 280046 61218 280102
rect 61274 280046 61342 280102
rect 61398 280046 69878 280102
rect 69934 280046 70002 280102
rect 70058 280046 78970 280102
rect 79026 280046 79094 280102
rect 79150 280046 79218 280102
rect 79274 280046 79342 280102
rect 79398 280046 96970 280102
rect 97026 280046 97094 280102
rect 97150 280046 97218 280102
rect 97274 280046 97342 280102
rect 97398 280046 100598 280102
rect 100654 280046 100722 280102
rect 100778 280046 131318 280102
rect 131374 280046 131442 280102
rect 131498 280046 162038 280102
rect 162094 280046 162162 280102
rect 162218 280046 192758 280102
rect 192814 280046 192882 280102
rect 192938 280046 223478 280102
rect 223534 280046 223602 280102
rect 223658 280046 254198 280102
rect 254254 280046 254322 280102
rect 254378 280046 284918 280102
rect 284974 280046 285042 280102
rect 285098 280046 315638 280102
rect 315694 280046 315762 280102
rect 315818 280046 346358 280102
rect 346414 280046 346482 280102
rect 346538 280046 377078 280102
rect 377134 280046 377202 280102
rect 377258 280046 407798 280102
rect 407854 280046 407922 280102
rect 407978 280046 438518 280102
rect 438574 280046 438642 280102
rect 438698 280046 469238 280102
rect 469294 280046 469362 280102
rect 469418 280046 499958 280102
rect 500014 280046 500082 280102
rect 500138 280046 530678 280102
rect 530734 280046 530802 280102
rect 530858 280046 564970 280102
rect 565026 280046 565094 280102
rect 565150 280046 565218 280102
rect 565274 280046 565342 280102
rect 565398 280046 582970 280102
rect 583026 280046 583094 280102
rect 583150 280046 583218 280102
rect 583274 280046 583342 280102
rect 583398 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect -1916 279978 597980 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 6970 279978
rect 7026 279922 7094 279978
rect 7150 279922 7218 279978
rect 7274 279922 7342 279978
rect 7398 279922 24970 279978
rect 25026 279922 25094 279978
rect 25150 279922 25218 279978
rect 25274 279922 25342 279978
rect 25398 279922 42970 279978
rect 43026 279922 43094 279978
rect 43150 279922 43218 279978
rect 43274 279922 43342 279978
rect 43398 279922 60970 279978
rect 61026 279922 61094 279978
rect 61150 279922 61218 279978
rect 61274 279922 61342 279978
rect 61398 279922 69878 279978
rect 69934 279922 70002 279978
rect 70058 279922 78970 279978
rect 79026 279922 79094 279978
rect 79150 279922 79218 279978
rect 79274 279922 79342 279978
rect 79398 279922 96970 279978
rect 97026 279922 97094 279978
rect 97150 279922 97218 279978
rect 97274 279922 97342 279978
rect 97398 279922 100598 279978
rect 100654 279922 100722 279978
rect 100778 279922 131318 279978
rect 131374 279922 131442 279978
rect 131498 279922 162038 279978
rect 162094 279922 162162 279978
rect 162218 279922 192758 279978
rect 192814 279922 192882 279978
rect 192938 279922 223478 279978
rect 223534 279922 223602 279978
rect 223658 279922 254198 279978
rect 254254 279922 254322 279978
rect 254378 279922 284918 279978
rect 284974 279922 285042 279978
rect 285098 279922 315638 279978
rect 315694 279922 315762 279978
rect 315818 279922 346358 279978
rect 346414 279922 346482 279978
rect 346538 279922 377078 279978
rect 377134 279922 377202 279978
rect 377258 279922 407798 279978
rect 407854 279922 407922 279978
rect 407978 279922 438518 279978
rect 438574 279922 438642 279978
rect 438698 279922 469238 279978
rect 469294 279922 469362 279978
rect 469418 279922 499958 279978
rect 500014 279922 500082 279978
rect 500138 279922 530678 279978
rect 530734 279922 530802 279978
rect 530858 279922 564970 279978
rect 565026 279922 565094 279978
rect 565150 279922 565218 279978
rect 565274 279922 565342 279978
rect 565398 279922 582970 279978
rect 583026 279922 583094 279978
rect 583150 279922 583218 279978
rect 583274 279922 583342 279978
rect 583398 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect -1916 279826 597980 279922
rect -1916 274350 597980 274446
rect -1916 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 3250 274350
rect 3306 274294 3374 274350
rect 3430 274294 3498 274350
rect 3554 274294 3622 274350
rect 3678 274294 21250 274350
rect 21306 274294 21374 274350
rect 21430 274294 21498 274350
rect 21554 274294 21622 274350
rect 21678 274294 39250 274350
rect 39306 274294 39374 274350
rect 39430 274294 39498 274350
rect 39554 274294 39622 274350
rect 39678 274294 54518 274350
rect 54574 274294 54642 274350
rect 54698 274294 57250 274350
rect 57306 274294 57374 274350
rect 57430 274294 57498 274350
rect 57554 274294 57622 274350
rect 57678 274294 75250 274350
rect 75306 274294 75374 274350
rect 75430 274294 75498 274350
rect 75554 274294 75622 274350
rect 75678 274294 85238 274350
rect 85294 274294 85362 274350
rect 85418 274294 93250 274350
rect 93306 274294 93374 274350
rect 93430 274294 93498 274350
rect 93554 274294 93622 274350
rect 93678 274294 111250 274350
rect 111306 274294 111374 274350
rect 111430 274294 111498 274350
rect 111554 274294 111622 274350
rect 111678 274294 115958 274350
rect 116014 274294 116082 274350
rect 116138 274294 146678 274350
rect 146734 274294 146802 274350
rect 146858 274294 177398 274350
rect 177454 274294 177522 274350
rect 177578 274294 208118 274350
rect 208174 274294 208242 274350
rect 208298 274294 238838 274350
rect 238894 274294 238962 274350
rect 239018 274294 269558 274350
rect 269614 274294 269682 274350
rect 269738 274294 300278 274350
rect 300334 274294 300402 274350
rect 300458 274294 330998 274350
rect 331054 274294 331122 274350
rect 331178 274294 361718 274350
rect 361774 274294 361842 274350
rect 361898 274294 392438 274350
rect 392494 274294 392562 274350
rect 392618 274294 423158 274350
rect 423214 274294 423282 274350
rect 423338 274294 453878 274350
rect 453934 274294 454002 274350
rect 454058 274294 484598 274350
rect 484654 274294 484722 274350
rect 484778 274294 515318 274350
rect 515374 274294 515442 274350
rect 515498 274294 546038 274350
rect 546094 274294 546162 274350
rect 546218 274294 561250 274350
rect 561306 274294 561374 274350
rect 561430 274294 561498 274350
rect 561554 274294 561622 274350
rect 561678 274294 579250 274350
rect 579306 274294 579374 274350
rect 579430 274294 579498 274350
rect 579554 274294 579622 274350
rect 579678 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597980 274350
rect -1916 274226 597980 274294
rect -1916 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 3250 274226
rect 3306 274170 3374 274226
rect 3430 274170 3498 274226
rect 3554 274170 3622 274226
rect 3678 274170 21250 274226
rect 21306 274170 21374 274226
rect 21430 274170 21498 274226
rect 21554 274170 21622 274226
rect 21678 274170 39250 274226
rect 39306 274170 39374 274226
rect 39430 274170 39498 274226
rect 39554 274170 39622 274226
rect 39678 274170 54518 274226
rect 54574 274170 54642 274226
rect 54698 274170 57250 274226
rect 57306 274170 57374 274226
rect 57430 274170 57498 274226
rect 57554 274170 57622 274226
rect 57678 274170 75250 274226
rect 75306 274170 75374 274226
rect 75430 274170 75498 274226
rect 75554 274170 75622 274226
rect 75678 274170 85238 274226
rect 85294 274170 85362 274226
rect 85418 274170 93250 274226
rect 93306 274170 93374 274226
rect 93430 274170 93498 274226
rect 93554 274170 93622 274226
rect 93678 274170 111250 274226
rect 111306 274170 111374 274226
rect 111430 274170 111498 274226
rect 111554 274170 111622 274226
rect 111678 274170 115958 274226
rect 116014 274170 116082 274226
rect 116138 274170 146678 274226
rect 146734 274170 146802 274226
rect 146858 274170 177398 274226
rect 177454 274170 177522 274226
rect 177578 274170 208118 274226
rect 208174 274170 208242 274226
rect 208298 274170 238838 274226
rect 238894 274170 238962 274226
rect 239018 274170 269558 274226
rect 269614 274170 269682 274226
rect 269738 274170 300278 274226
rect 300334 274170 300402 274226
rect 300458 274170 330998 274226
rect 331054 274170 331122 274226
rect 331178 274170 361718 274226
rect 361774 274170 361842 274226
rect 361898 274170 392438 274226
rect 392494 274170 392562 274226
rect 392618 274170 423158 274226
rect 423214 274170 423282 274226
rect 423338 274170 453878 274226
rect 453934 274170 454002 274226
rect 454058 274170 484598 274226
rect 484654 274170 484722 274226
rect 484778 274170 515318 274226
rect 515374 274170 515442 274226
rect 515498 274170 546038 274226
rect 546094 274170 546162 274226
rect 546218 274170 561250 274226
rect 561306 274170 561374 274226
rect 561430 274170 561498 274226
rect 561554 274170 561622 274226
rect 561678 274170 579250 274226
rect 579306 274170 579374 274226
rect 579430 274170 579498 274226
rect 579554 274170 579622 274226
rect 579678 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597980 274226
rect -1916 274102 597980 274170
rect -1916 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 3250 274102
rect 3306 274046 3374 274102
rect 3430 274046 3498 274102
rect 3554 274046 3622 274102
rect 3678 274046 21250 274102
rect 21306 274046 21374 274102
rect 21430 274046 21498 274102
rect 21554 274046 21622 274102
rect 21678 274046 39250 274102
rect 39306 274046 39374 274102
rect 39430 274046 39498 274102
rect 39554 274046 39622 274102
rect 39678 274046 54518 274102
rect 54574 274046 54642 274102
rect 54698 274046 57250 274102
rect 57306 274046 57374 274102
rect 57430 274046 57498 274102
rect 57554 274046 57622 274102
rect 57678 274046 75250 274102
rect 75306 274046 75374 274102
rect 75430 274046 75498 274102
rect 75554 274046 75622 274102
rect 75678 274046 85238 274102
rect 85294 274046 85362 274102
rect 85418 274046 93250 274102
rect 93306 274046 93374 274102
rect 93430 274046 93498 274102
rect 93554 274046 93622 274102
rect 93678 274046 111250 274102
rect 111306 274046 111374 274102
rect 111430 274046 111498 274102
rect 111554 274046 111622 274102
rect 111678 274046 115958 274102
rect 116014 274046 116082 274102
rect 116138 274046 146678 274102
rect 146734 274046 146802 274102
rect 146858 274046 177398 274102
rect 177454 274046 177522 274102
rect 177578 274046 208118 274102
rect 208174 274046 208242 274102
rect 208298 274046 238838 274102
rect 238894 274046 238962 274102
rect 239018 274046 269558 274102
rect 269614 274046 269682 274102
rect 269738 274046 300278 274102
rect 300334 274046 300402 274102
rect 300458 274046 330998 274102
rect 331054 274046 331122 274102
rect 331178 274046 361718 274102
rect 361774 274046 361842 274102
rect 361898 274046 392438 274102
rect 392494 274046 392562 274102
rect 392618 274046 423158 274102
rect 423214 274046 423282 274102
rect 423338 274046 453878 274102
rect 453934 274046 454002 274102
rect 454058 274046 484598 274102
rect 484654 274046 484722 274102
rect 484778 274046 515318 274102
rect 515374 274046 515442 274102
rect 515498 274046 546038 274102
rect 546094 274046 546162 274102
rect 546218 274046 561250 274102
rect 561306 274046 561374 274102
rect 561430 274046 561498 274102
rect 561554 274046 561622 274102
rect 561678 274046 579250 274102
rect 579306 274046 579374 274102
rect 579430 274046 579498 274102
rect 579554 274046 579622 274102
rect 579678 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597980 274102
rect -1916 273978 597980 274046
rect -1916 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 3250 273978
rect 3306 273922 3374 273978
rect 3430 273922 3498 273978
rect 3554 273922 3622 273978
rect 3678 273922 21250 273978
rect 21306 273922 21374 273978
rect 21430 273922 21498 273978
rect 21554 273922 21622 273978
rect 21678 273922 39250 273978
rect 39306 273922 39374 273978
rect 39430 273922 39498 273978
rect 39554 273922 39622 273978
rect 39678 273922 54518 273978
rect 54574 273922 54642 273978
rect 54698 273922 57250 273978
rect 57306 273922 57374 273978
rect 57430 273922 57498 273978
rect 57554 273922 57622 273978
rect 57678 273922 75250 273978
rect 75306 273922 75374 273978
rect 75430 273922 75498 273978
rect 75554 273922 75622 273978
rect 75678 273922 85238 273978
rect 85294 273922 85362 273978
rect 85418 273922 93250 273978
rect 93306 273922 93374 273978
rect 93430 273922 93498 273978
rect 93554 273922 93622 273978
rect 93678 273922 111250 273978
rect 111306 273922 111374 273978
rect 111430 273922 111498 273978
rect 111554 273922 111622 273978
rect 111678 273922 115958 273978
rect 116014 273922 116082 273978
rect 116138 273922 146678 273978
rect 146734 273922 146802 273978
rect 146858 273922 177398 273978
rect 177454 273922 177522 273978
rect 177578 273922 208118 273978
rect 208174 273922 208242 273978
rect 208298 273922 238838 273978
rect 238894 273922 238962 273978
rect 239018 273922 269558 273978
rect 269614 273922 269682 273978
rect 269738 273922 300278 273978
rect 300334 273922 300402 273978
rect 300458 273922 330998 273978
rect 331054 273922 331122 273978
rect 331178 273922 361718 273978
rect 361774 273922 361842 273978
rect 361898 273922 392438 273978
rect 392494 273922 392562 273978
rect 392618 273922 423158 273978
rect 423214 273922 423282 273978
rect 423338 273922 453878 273978
rect 453934 273922 454002 273978
rect 454058 273922 484598 273978
rect 484654 273922 484722 273978
rect 484778 273922 515318 273978
rect 515374 273922 515442 273978
rect 515498 273922 546038 273978
rect 546094 273922 546162 273978
rect 546218 273922 561250 273978
rect 561306 273922 561374 273978
rect 561430 273922 561498 273978
rect 561554 273922 561622 273978
rect 561678 273922 579250 273978
rect 579306 273922 579374 273978
rect 579430 273922 579498 273978
rect 579554 273922 579622 273978
rect 579678 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597980 273978
rect -1916 273826 597980 273922
rect -1916 262350 597980 262446
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 6970 262350
rect 7026 262294 7094 262350
rect 7150 262294 7218 262350
rect 7274 262294 7342 262350
rect 7398 262294 24970 262350
rect 25026 262294 25094 262350
rect 25150 262294 25218 262350
rect 25274 262294 25342 262350
rect 25398 262294 42970 262350
rect 43026 262294 43094 262350
rect 43150 262294 43218 262350
rect 43274 262294 43342 262350
rect 43398 262294 60970 262350
rect 61026 262294 61094 262350
rect 61150 262294 61218 262350
rect 61274 262294 61342 262350
rect 61398 262294 69878 262350
rect 69934 262294 70002 262350
rect 70058 262294 78970 262350
rect 79026 262294 79094 262350
rect 79150 262294 79218 262350
rect 79274 262294 79342 262350
rect 79398 262294 96970 262350
rect 97026 262294 97094 262350
rect 97150 262294 97218 262350
rect 97274 262294 97342 262350
rect 97398 262294 100598 262350
rect 100654 262294 100722 262350
rect 100778 262294 131318 262350
rect 131374 262294 131442 262350
rect 131498 262294 162038 262350
rect 162094 262294 162162 262350
rect 162218 262294 192758 262350
rect 192814 262294 192882 262350
rect 192938 262294 223478 262350
rect 223534 262294 223602 262350
rect 223658 262294 254198 262350
rect 254254 262294 254322 262350
rect 254378 262294 284918 262350
rect 284974 262294 285042 262350
rect 285098 262294 315638 262350
rect 315694 262294 315762 262350
rect 315818 262294 346358 262350
rect 346414 262294 346482 262350
rect 346538 262294 377078 262350
rect 377134 262294 377202 262350
rect 377258 262294 407798 262350
rect 407854 262294 407922 262350
rect 407978 262294 438518 262350
rect 438574 262294 438642 262350
rect 438698 262294 469238 262350
rect 469294 262294 469362 262350
rect 469418 262294 499958 262350
rect 500014 262294 500082 262350
rect 500138 262294 530678 262350
rect 530734 262294 530802 262350
rect 530858 262294 564970 262350
rect 565026 262294 565094 262350
rect 565150 262294 565218 262350
rect 565274 262294 565342 262350
rect 565398 262294 582970 262350
rect 583026 262294 583094 262350
rect 583150 262294 583218 262350
rect 583274 262294 583342 262350
rect 583398 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect -1916 262226 597980 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 6970 262226
rect 7026 262170 7094 262226
rect 7150 262170 7218 262226
rect 7274 262170 7342 262226
rect 7398 262170 24970 262226
rect 25026 262170 25094 262226
rect 25150 262170 25218 262226
rect 25274 262170 25342 262226
rect 25398 262170 42970 262226
rect 43026 262170 43094 262226
rect 43150 262170 43218 262226
rect 43274 262170 43342 262226
rect 43398 262170 60970 262226
rect 61026 262170 61094 262226
rect 61150 262170 61218 262226
rect 61274 262170 61342 262226
rect 61398 262170 69878 262226
rect 69934 262170 70002 262226
rect 70058 262170 78970 262226
rect 79026 262170 79094 262226
rect 79150 262170 79218 262226
rect 79274 262170 79342 262226
rect 79398 262170 96970 262226
rect 97026 262170 97094 262226
rect 97150 262170 97218 262226
rect 97274 262170 97342 262226
rect 97398 262170 100598 262226
rect 100654 262170 100722 262226
rect 100778 262170 131318 262226
rect 131374 262170 131442 262226
rect 131498 262170 162038 262226
rect 162094 262170 162162 262226
rect 162218 262170 192758 262226
rect 192814 262170 192882 262226
rect 192938 262170 223478 262226
rect 223534 262170 223602 262226
rect 223658 262170 254198 262226
rect 254254 262170 254322 262226
rect 254378 262170 284918 262226
rect 284974 262170 285042 262226
rect 285098 262170 315638 262226
rect 315694 262170 315762 262226
rect 315818 262170 346358 262226
rect 346414 262170 346482 262226
rect 346538 262170 377078 262226
rect 377134 262170 377202 262226
rect 377258 262170 407798 262226
rect 407854 262170 407922 262226
rect 407978 262170 438518 262226
rect 438574 262170 438642 262226
rect 438698 262170 469238 262226
rect 469294 262170 469362 262226
rect 469418 262170 499958 262226
rect 500014 262170 500082 262226
rect 500138 262170 530678 262226
rect 530734 262170 530802 262226
rect 530858 262170 564970 262226
rect 565026 262170 565094 262226
rect 565150 262170 565218 262226
rect 565274 262170 565342 262226
rect 565398 262170 582970 262226
rect 583026 262170 583094 262226
rect 583150 262170 583218 262226
rect 583274 262170 583342 262226
rect 583398 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect -1916 262102 597980 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 6970 262102
rect 7026 262046 7094 262102
rect 7150 262046 7218 262102
rect 7274 262046 7342 262102
rect 7398 262046 24970 262102
rect 25026 262046 25094 262102
rect 25150 262046 25218 262102
rect 25274 262046 25342 262102
rect 25398 262046 42970 262102
rect 43026 262046 43094 262102
rect 43150 262046 43218 262102
rect 43274 262046 43342 262102
rect 43398 262046 60970 262102
rect 61026 262046 61094 262102
rect 61150 262046 61218 262102
rect 61274 262046 61342 262102
rect 61398 262046 69878 262102
rect 69934 262046 70002 262102
rect 70058 262046 78970 262102
rect 79026 262046 79094 262102
rect 79150 262046 79218 262102
rect 79274 262046 79342 262102
rect 79398 262046 96970 262102
rect 97026 262046 97094 262102
rect 97150 262046 97218 262102
rect 97274 262046 97342 262102
rect 97398 262046 100598 262102
rect 100654 262046 100722 262102
rect 100778 262046 131318 262102
rect 131374 262046 131442 262102
rect 131498 262046 162038 262102
rect 162094 262046 162162 262102
rect 162218 262046 192758 262102
rect 192814 262046 192882 262102
rect 192938 262046 223478 262102
rect 223534 262046 223602 262102
rect 223658 262046 254198 262102
rect 254254 262046 254322 262102
rect 254378 262046 284918 262102
rect 284974 262046 285042 262102
rect 285098 262046 315638 262102
rect 315694 262046 315762 262102
rect 315818 262046 346358 262102
rect 346414 262046 346482 262102
rect 346538 262046 377078 262102
rect 377134 262046 377202 262102
rect 377258 262046 407798 262102
rect 407854 262046 407922 262102
rect 407978 262046 438518 262102
rect 438574 262046 438642 262102
rect 438698 262046 469238 262102
rect 469294 262046 469362 262102
rect 469418 262046 499958 262102
rect 500014 262046 500082 262102
rect 500138 262046 530678 262102
rect 530734 262046 530802 262102
rect 530858 262046 564970 262102
rect 565026 262046 565094 262102
rect 565150 262046 565218 262102
rect 565274 262046 565342 262102
rect 565398 262046 582970 262102
rect 583026 262046 583094 262102
rect 583150 262046 583218 262102
rect 583274 262046 583342 262102
rect 583398 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect -1916 261978 597980 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 6970 261978
rect 7026 261922 7094 261978
rect 7150 261922 7218 261978
rect 7274 261922 7342 261978
rect 7398 261922 24970 261978
rect 25026 261922 25094 261978
rect 25150 261922 25218 261978
rect 25274 261922 25342 261978
rect 25398 261922 42970 261978
rect 43026 261922 43094 261978
rect 43150 261922 43218 261978
rect 43274 261922 43342 261978
rect 43398 261922 60970 261978
rect 61026 261922 61094 261978
rect 61150 261922 61218 261978
rect 61274 261922 61342 261978
rect 61398 261922 69878 261978
rect 69934 261922 70002 261978
rect 70058 261922 78970 261978
rect 79026 261922 79094 261978
rect 79150 261922 79218 261978
rect 79274 261922 79342 261978
rect 79398 261922 96970 261978
rect 97026 261922 97094 261978
rect 97150 261922 97218 261978
rect 97274 261922 97342 261978
rect 97398 261922 100598 261978
rect 100654 261922 100722 261978
rect 100778 261922 131318 261978
rect 131374 261922 131442 261978
rect 131498 261922 162038 261978
rect 162094 261922 162162 261978
rect 162218 261922 192758 261978
rect 192814 261922 192882 261978
rect 192938 261922 223478 261978
rect 223534 261922 223602 261978
rect 223658 261922 254198 261978
rect 254254 261922 254322 261978
rect 254378 261922 284918 261978
rect 284974 261922 285042 261978
rect 285098 261922 315638 261978
rect 315694 261922 315762 261978
rect 315818 261922 346358 261978
rect 346414 261922 346482 261978
rect 346538 261922 377078 261978
rect 377134 261922 377202 261978
rect 377258 261922 407798 261978
rect 407854 261922 407922 261978
rect 407978 261922 438518 261978
rect 438574 261922 438642 261978
rect 438698 261922 469238 261978
rect 469294 261922 469362 261978
rect 469418 261922 499958 261978
rect 500014 261922 500082 261978
rect 500138 261922 530678 261978
rect 530734 261922 530802 261978
rect 530858 261922 564970 261978
rect 565026 261922 565094 261978
rect 565150 261922 565218 261978
rect 565274 261922 565342 261978
rect 565398 261922 582970 261978
rect 583026 261922 583094 261978
rect 583150 261922 583218 261978
rect 583274 261922 583342 261978
rect 583398 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect -1916 261826 597980 261922
rect -1916 256350 597980 256446
rect -1916 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 3250 256350
rect 3306 256294 3374 256350
rect 3430 256294 3498 256350
rect 3554 256294 3622 256350
rect 3678 256294 21250 256350
rect 21306 256294 21374 256350
rect 21430 256294 21498 256350
rect 21554 256294 21622 256350
rect 21678 256294 39250 256350
rect 39306 256294 39374 256350
rect 39430 256294 39498 256350
rect 39554 256294 39622 256350
rect 39678 256294 54518 256350
rect 54574 256294 54642 256350
rect 54698 256294 57250 256350
rect 57306 256294 57374 256350
rect 57430 256294 57498 256350
rect 57554 256294 57622 256350
rect 57678 256294 75250 256350
rect 75306 256294 75374 256350
rect 75430 256294 75498 256350
rect 75554 256294 75622 256350
rect 75678 256294 85238 256350
rect 85294 256294 85362 256350
rect 85418 256294 93250 256350
rect 93306 256294 93374 256350
rect 93430 256294 93498 256350
rect 93554 256294 93622 256350
rect 93678 256294 111250 256350
rect 111306 256294 111374 256350
rect 111430 256294 111498 256350
rect 111554 256294 111622 256350
rect 111678 256294 115958 256350
rect 116014 256294 116082 256350
rect 116138 256294 146678 256350
rect 146734 256294 146802 256350
rect 146858 256294 177398 256350
rect 177454 256294 177522 256350
rect 177578 256294 208118 256350
rect 208174 256294 208242 256350
rect 208298 256294 238838 256350
rect 238894 256294 238962 256350
rect 239018 256294 269558 256350
rect 269614 256294 269682 256350
rect 269738 256294 300278 256350
rect 300334 256294 300402 256350
rect 300458 256294 330998 256350
rect 331054 256294 331122 256350
rect 331178 256294 361718 256350
rect 361774 256294 361842 256350
rect 361898 256294 392438 256350
rect 392494 256294 392562 256350
rect 392618 256294 423158 256350
rect 423214 256294 423282 256350
rect 423338 256294 453878 256350
rect 453934 256294 454002 256350
rect 454058 256294 484598 256350
rect 484654 256294 484722 256350
rect 484778 256294 515318 256350
rect 515374 256294 515442 256350
rect 515498 256294 546038 256350
rect 546094 256294 546162 256350
rect 546218 256294 561250 256350
rect 561306 256294 561374 256350
rect 561430 256294 561498 256350
rect 561554 256294 561622 256350
rect 561678 256294 579250 256350
rect 579306 256294 579374 256350
rect 579430 256294 579498 256350
rect 579554 256294 579622 256350
rect 579678 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597980 256350
rect -1916 256226 597980 256294
rect -1916 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 3250 256226
rect 3306 256170 3374 256226
rect 3430 256170 3498 256226
rect 3554 256170 3622 256226
rect 3678 256170 21250 256226
rect 21306 256170 21374 256226
rect 21430 256170 21498 256226
rect 21554 256170 21622 256226
rect 21678 256170 39250 256226
rect 39306 256170 39374 256226
rect 39430 256170 39498 256226
rect 39554 256170 39622 256226
rect 39678 256170 54518 256226
rect 54574 256170 54642 256226
rect 54698 256170 57250 256226
rect 57306 256170 57374 256226
rect 57430 256170 57498 256226
rect 57554 256170 57622 256226
rect 57678 256170 75250 256226
rect 75306 256170 75374 256226
rect 75430 256170 75498 256226
rect 75554 256170 75622 256226
rect 75678 256170 85238 256226
rect 85294 256170 85362 256226
rect 85418 256170 93250 256226
rect 93306 256170 93374 256226
rect 93430 256170 93498 256226
rect 93554 256170 93622 256226
rect 93678 256170 111250 256226
rect 111306 256170 111374 256226
rect 111430 256170 111498 256226
rect 111554 256170 111622 256226
rect 111678 256170 115958 256226
rect 116014 256170 116082 256226
rect 116138 256170 146678 256226
rect 146734 256170 146802 256226
rect 146858 256170 177398 256226
rect 177454 256170 177522 256226
rect 177578 256170 208118 256226
rect 208174 256170 208242 256226
rect 208298 256170 238838 256226
rect 238894 256170 238962 256226
rect 239018 256170 269558 256226
rect 269614 256170 269682 256226
rect 269738 256170 300278 256226
rect 300334 256170 300402 256226
rect 300458 256170 330998 256226
rect 331054 256170 331122 256226
rect 331178 256170 361718 256226
rect 361774 256170 361842 256226
rect 361898 256170 392438 256226
rect 392494 256170 392562 256226
rect 392618 256170 423158 256226
rect 423214 256170 423282 256226
rect 423338 256170 453878 256226
rect 453934 256170 454002 256226
rect 454058 256170 484598 256226
rect 484654 256170 484722 256226
rect 484778 256170 515318 256226
rect 515374 256170 515442 256226
rect 515498 256170 546038 256226
rect 546094 256170 546162 256226
rect 546218 256170 561250 256226
rect 561306 256170 561374 256226
rect 561430 256170 561498 256226
rect 561554 256170 561622 256226
rect 561678 256170 579250 256226
rect 579306 256170 579374 256226
rect 579430 256170 579498 256226
rect 579554 256170 579622 256226
rect 579678 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597980 256226
rect -1916 256102 597980 256170
rect -1916 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 3250 256102
rect 3306 256046 3374 256102
rect 3430 256046 3498 256102
rect 3554 256046 3622 256102
rect 3678 256046 21250 256102
rect 21306 256046 21374 256102
rect 21430 256046 21498 256102
rect 21554 256046 21622 256102
rect 21678 256046 39250 256102
rect 39306 256046 39374 256102
rect 39430 256046 39498 256102
rect 39554 256046 39622 256102
rect 39678 256046 54518 256102
rect 54574 256046 54642 256102
rect 54698 256046 57250 256102
rect 57306 256046 57374 256102
rect 57430 256046 57498 256102
rect 57554 256046 57622 256102
rect 57678 256046 75250 256102
rect 75306 256046 75374 256102
rect 75430 256046 75498 256102
rect 75554 256046 75622 256102
rect 75678 256046 85238 256102
rect 85294 256046 85362 256102
rect 85418 256046 93250 256102
rect 93306 256046 93374 256102
rect 93430 256046 93498 256102
rect 93554 256046 93622 256102
rect 93678 256046 111250 256102
rect 111306 256046 111374 256102
rect 111430 256046 111498 256102
rect 111554 256046 111622 256102
rect 111678 256046 115958 256102
rect 116014 256046 116082 256102
rect 116138 256046 146678 256102
rect 146734 256046 146802 256102
rect 146858 256046 177398 256102
rect 177454 256046 177522 256102
rect 177578 256046 208118 256102
rect 208174 256046 208242 256102
rect 208298 256046 238838 256102
rect 238894 256046 238962 256102
rect 239018 256046 269558 256102
rect 269614 256046 269682 256102
rect 269738 256046 300278 256102
rect 300334 256046 300402 256102
rect 300458 256046 330998 256102
rect 331054 256046 331122 256102
rect 331178 256046 361718 256102
rect 361774 256046 361842 256102
rect 361898 256046 392438 256102
rect 392494 256046 392562 256102
rect 392618 256046 423158 256102
rect 423214 256046 423282 256102
rect 423338 256046 453878 256102
rect 453934 256046 454002 256102
rect 454058 256046 484598 256102
rect 484654 256046 484722 256102
rect 484778 256046 515318 256102
rect 515374 256046 515442 256102
rect 515498 256046 546038 256102
rect 546094 256046 546162 256102
rect 546218 256046 561250 256102
rect 561306 256046 561374 256102
rect 561430 256046 561498 256102
rect 561554 256046 561622 256102
rect 561678 256046 579250 256102
rect 579306 256046 579374 256102
rect 579430 256046 579498 256102
rect 579554 256046 579622 256102
rect 579678 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597980 256102
rect -1916 255978 597980 256046
rect -1916 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 3250 255978
rect 3306 255922 3374 255978
rect 3430 255922 3498 255978
rect 3554 255922 3622 255978
rect 3678 255922 21250 255978
rect 21306 255922 21374 255978
rect 21430 255922 21498 255978
rect 21554 255922 21622 255978
rect 21678 255922 39250 255978
rect 39306 255922 39374 255978
rect 39430 255922 39498 255978
rect 39554 255922 39622 255978
rect 39678 255922 54518 255978
rect 54574 255922 54642 255978
rect 54698 255922 57250 255978
rect 57306 255922 57374 255978
rect 57430 255922 57498 255978
rect 57554 255922 57622 255978
rect 57678 255922 75250 255978
rect 75306 255922 75374 255978
rect 75430 255922 75498 255978
rect 75554 255922 75622 255978
rect 75678 255922 85238 255978
rect 85294 255922 85362 255978
rect 85418 255922 93250 255978
rect 93306 255922 93374 255978
rect 93430 255922 93498 255978
rect 93554 255922 93622 255978
rect 93678 255922 111250 255978
rect 111306 255922 111374 255978
rect 111430 255922 111498 255978
rect 111554 255922 111622 255978
rect 111678 255922 115958 255978
rect 116014 255922 116082 255978
rect 116138 255922 146678 255978
rect 146734 255922 146802 255978
rect 146858 255922 177398 255978
rect 177454 255922 177522 255978
rect 177578 255922 208118 255978
rect 208174 255922 208242 255978
rect 208298 255922 238838 255978
rect 238894 255922 238962 255978
rect 239018 255922 269558 255978
rect 269614 255922 269682 255978
rect 269738 255922 300278 255978
rect 300334 255922 300402 255978
rect 300458 255922 330998 255978
rect 331054 255922 331122 255978
rect 331178 255922 361718 255978
rect 361774 255922 361842 255978
rect 361898 255922 392438 255978
rect 392494 255922 392562 255978
rect 392618 255922 423158 255978
rect 423214 255922 423282 255978
rect 423338 255922 453878 255978
rect 453934 255922 454002 255978
rect 454058 255922 484598 255978
rect 484654 255922 484722 255978
rect 484778 255922 515318 255978
rect 515374 255922 515442 255978
rect 515498 255922 546038 255978
rect 546094 255922 546162 255978
rect 546218 255922 561250 255978
rect 561306 255922 561374 255978
rect 561430 255922 561498 255978
rect 561554 255922 561622 255978
rect 561678 255922 579250 255978
rect 579306 255922 579374 255978
rect 579430 255922 579498 255978
rect 579554 255922 579622 255978
rect 579678 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597980 255978
rect -1916 255826 597980 255922
rect -1916 244350 597980 244446
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 6970 244350
rect 7026 244294 7094 244350
rect 7150 244294 7218 244350
rect 7274 244294 7342 244350
rect 7398 244294 24970 244350
rect 25026 244294 25094 244350
rect 25150 244294 25218 244350
rect 25274 244294 25342 244350
rect 25398 244294 42970 244350
rect 43026 244294 43094 244350
rect 43150 244294 43218 244350
rect 43274 244294 43342 244350
rect 43398 244294 60970 244350
rect 61026 244294 61094 244350
rect 61150 244294 61218 244350
rect 61274 244294 61342 244350
rect 61398 244294 69878 244350
rect 69934 244294 70002 244350
rect 70058 244294 78970 244350
rect 79026 244294 79094 244350
rect 79150 244294 79218 244350
rect 79274 244294 79342 244350
rect 79398 244294 96970 244350
rect 97026 244294 97094 244350
rect 97150 244294 97218 244350
rect 97274 244294 97342 244350
rect 97398 244294 100598 244350
rect 100654 244294 100722 244350
rect 100778 244294 131318 244350
rect 131374 244294 131442 244350
rect 131498 244294 162038 244350
rect 162094 244294 162162 244350
rect 162218 244294 192758 244350
rect 192814 244294 192882 244350
rect 192938 244294 223478 244350
rect 223534 244294 223602 244350
rect 223658 244294 254198 244350
rect 254254 244294 254322 244350
rect 254378 244294 284918 244350
rect 284974 244294 285042 244350
rect 285098 244294 315638 244350
rect 315694 244294 315762 244350
rect 315818 244294 346358 244350
rect 346414 244294 346482 244350
rect 346538 244294 377078 244350
rect 377134 244294 377202 244350
rect 377258 244294 407798 244350
rect 407854 244294 407922 244350
rect 407978 244294 438518 244350
rect 438574 244294 438642 244350
rect 438698 244294 469238 244350
rect 469294 244294 469362 244350
rect 469418 244294 499958 244350
rect 500014 244294 500082 244350
rect 500138 244294 530678 244350
rect 530734 244294 530802 244350
rect 530858 244294 564970 244350
rect 565026 244294 565094 244350
rect 565150 244294 565218 244350
rect 565274 244294 565342 244350
rect 565398 244294 582970 244350
rect 583026 244294 583094 244350
rect 583150 244294 583218 244350
rect 583274 244294 583342 244350
rect 583398 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect -1916 244226 597980 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 6970 244226
rect 7026 244170 7094 244226
rect 7150 244170 7218 244226
rect 7274 244170 7342 244226
rect 7398 244170 24970 244226
rect 25026 244170 25094 244226
rect 25150 244170 25218 244226
rect 25274 244170 25342 244226
rect 25398 244170 42970 244226
rect 43026 244170 43094 244226
rect 43150 244170 43218 244226
rect 43274 244170 43342 244226
rect 43398 244170 60970 244226
rect 61026 244170 61094 244226
rect 61150 244170 61218 244226
rect 61274 244170 61342 244226
rect 61398 244170 69878 244226
rect 69934 244170 70002 244226
rect 70058 244170 78970 244226
rect 79026 244170 79094 244226
rect 79150 244170 79218 244226
rect 79274 244170 79342 244226
rect 79398 244170 96970 244226
rect 97026 244170 97094 244226
rect 97150 244170 97218 244226
rect 97274 244170 97342 244226
rect 97398 244170 100598 244226
rect 100654 244170 100722 244226
rect 100778 244170 131318 244226
rect 131374 244170 131442 244226
rect 131498 244170 162038 244226
rect 162094 244170 162162 244226
rect 162218 244170 192758 244226
rect 192814 244170 192882 244226
rect 192938 244170 223478 244226
rect 223534 244170 223602 244226
rect 223658 244170 254198 244226
rect 254254 244170 254322 244226
rect 254378 244170 284918 244226
rect 284974 244170 285042 244226
rect 285098 244170 315638 244226
rect 315694 244170 315762 244226
rect 315818 244170 346358 244226
rect 346414 244170 346482 244226
rect 346538 244170 377078 244226
rect 377134 244170 377202 244226
rect 377258 244170 407798 244226
rect 407854 244170 407922 244226
rect 407978 244170 438518 244226
rect 438574 244170 438642 244226
rect 438698 244170 469238 244226
rect 469294 244170 469362 244226
rect 469418 244170 499958 244226
rect 500014 244170 500082 244226
rect 500138 244170 530678 244226
rect 530734 244170 530802 244226
rect 530858 244170 564970 244226
rect 565026 244170 565094 244226
rect 565150 244170 565218 244226
rect 565274 244170 565342 244226
rect 565398 244170 582970 244226
rect 583026 244170 583094 244226
rect 583150 244170 583218 244226
rect 583274 244170 583342 244226
rect 583398 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect -1916 244102 597980 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 6970 244102
rect 7026 244046 7094 244102
rect 7150 244046 7218 244102
rect 7274 244046 7342 244102
rect 7398 244046 24970 244102
rect 25026 244046 25094 244102
rect 25150 244046 25218 244102
rect 25274 244046 25342 244102
rect 25398 244046 42970 244102
rect 43026 244046 43094 244102
rect 43150 244046 43218 244102
rect 43274 244046 43342 244102
rect 43398 244046 60970 244102
rect 61026 244046 61094 244102
rect 61150 244046 61218 244102
rect 61274 244046 61342 244102
rect 61398 244046 69878 244102
rect 69934 244046 70002 244102
rect 70058 244046 78970 244102
rect 79026 244046 79094 244102
rect 79150 244046 79218 244102
rect 79274 244046 79342 244102
rect 79398 244046 96970 244102
rect 97026 244046 97094 244102
rect 97150 244046 97218 244102
rect 97274 244046 97342 244102
rect 97398 244046 100598 244102
rect 100654 244046 100722 244102
rect 100778 244046 131318 244102
rect 131374 244046 131442 244102
rect 131498 244046 162038 244102
rect 162094 244046 162162 244102
rect 162218 244046 192758 244102
rect 192814 244046 192882 244102
rect 192938 244046 223478 244102
rect 223534 244046 223602 244102
rect 223658 244046 254198 244102
rect 254254 244046 254322 244102
rect 254378 244046 284918 244102
rect 284974 244046 285042 244102
rect 285098 244046 315638 244102
rect 315694 244046 315762 244102
rect 315818 244046 346358 244102
rect 346414 244046 346482 244102
rect 346538 244046 377078 244102
rect 377134 244046 377202 244102
rect 377258 244046 407798 244102
rect 407854 244046 407922 244102
rect 407978 244046 438518 244102
rect 438574 244046 438642 244102
rect 438698 244046 469238 244102
rect 469294 244046 469362 244102
rect 469418 244046 499958 244102
rect 500014 244046 500082 244102
rect 500138 244046 530678 244102
rect 530734 244046 530802 244102
rect 530858 244046 564970 244102
rect 565026 244046 565094 244102
rect 565150 244046 565218 244102
rect 565274 244046 565342 244102
rect 565398 244046 582970 244102
rect 583026 244046 583094 244102
rect 583150 244046 583218 244102
rect 583274 244046 583342 244102
rect 583398 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect -1916 243978 597980 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 6970 243978
rect 7026 243922 7094 243978
rect 7150 243922 7218 243978
rect 7274 243922 7342 243978
rect 7398 243922 24970 243978
rect 25026 243922 25094 243978
rect 25150 243922 25218 243978
rect 25274 243922 25342 243978
rect 25398 243922 42970 243978
rect 43026 243922 43094 243978
rect 43150 243922 43218 243978
rect 43274 243922 43342 243978
rect 43398 243922 60970 243978
rect 61026 243922 61094 243978
rect 61150 243922 61218 243978
rect 61274 243922 61342 243978
rect 61398 243922 69878 243978
rect 69934 243922 70002 243978
rect 70058 243922 78970 243978
rect 79026 243922 79094 243978
rect 79150 243922 79218 243978
rect 79274 243922 79342 243978
rect 79398 243922 96970 243978
rect 97026 243922 97094 243978
rect 97150 243922 97218 243978
rect 97274 243922 97342 243978
rect 97398 243922 100598 243978
rect 100654 243922 100722 243978
rect 100778 243922 131318 243978
rect 131374 243922 131442 243978
rect 131498 243922 162038 243978
rect 162094 243922 162162 243978
rect 162218 243922 192758 243978
rect 192814 243922 192882 243978
rect 192938 243922 223478 243978
rect 223534 243922 223602 243978
rect 223658 243922 254198 243978
rect 254254 243922 254322 243978
rect 254378 243922 284918 243978
rect 284974 243922 285042 243978
rect 285098 243922 315638 243978
rect 315694 243922 315762 243978
rect 315818 243922 346358 243978
rect 346414 243922 346482 243978
rect 346538 243922 377078 243978
rect 377134 243922 377202 243978
rect 377258 243922 407798 243978
rect 407854 243922 407922 243978
rect 407978 243922 438518 243978
rect 438574 243922 438642 243978
rect 438698 243922 469238 243978
rect 469294 243922 469362 243978
rect 469418 243922 499958 243978
rect 500014 243922 500082 243978
rect 500138 243922 530678 243978
rect 530734 243922 530802 243978
rect 530858 243922 564970 243978
rect 565026 243922 565094 243978
rect 565150 243922 565218 243978
rect 565274 243922 565342 243978
rect 565398 243922 582970 243978
rect 583026 243922 583094 243978
rect 583150 243922 583218 243978
rect 583274 243922 583342 243978
rect 583398 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect -1916 243826 597980 243922
rect -1916 238350 597980 238446
rect -1916 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 3250 238350
rect 3306 238294 3374 238350
rect 3430 238294 3498 238350
rect 3554 238294 3622 238350
rect 3678 238294 21250 238350
rect 21306 238294 21374 238350
rect 21430 238294 21498 238350
rect 21554 238294 21622 238350
rect 21678 238294 39250 238350
rect 39306 238294 39374 238350
rect 39430 238294 39498 238350
rect 39554 238294 39622 238350
rect 39678 238294 54518 238350
rect 54574 238294 54642 238350
rect 54698 238294 57250 238350
rect 57306 238294 57374 238350
rect 57430 238294 57498 238350
rect 57554 238294 57622 238350
rect 57678 238294 75250 238350
rect 75306 238294 75374 238350
rect 75430 238294 75498 238350
rect 75554 238294 75622 238350
rect 75678 238294 85238 238350
rect 85294 238294 85362 238350
rect 85418 238294 93250 238350
rect 93306 238294 93374 238350
rect 93430 238294 93498 238350
rect 93554 238294 93622 238350
rect 93678 238294 111250 238350
rect 111306 238294 111374 238350
rect 111430 238294 111498 238350
rect 111554 238294 111622 238350
rect 111678 238294 115958 238350
rect 116014 238294 116082 238350
rect 116138 238294 146678 238350
rect 146734 238294 146802 238350
rect 146858 238294 177398 238350
rect 177454 238294 177522 238350
rect 177578 238294 208118 238350
rect 208174 238294 208242 238350
rect 208298 238294 238838 238350
rect 238894 238294 238962 238350
rect 239018 238294 269558 238350
rect 269614 238294 269682 238350
rect 269738 238294 300278 238350
rect 300334 238294 300402 238350
rect 300458 238294 330998 238350
rect 331054 238294 331122 238350
rect 331178 238294 361718 238350
rect 361774 238294 361842 238350
rect 361898 238294 392438 238350
rect 392494 238294 392562 238350
rect 392618 238294 423158 238350
rect 423214 238294 423282 238350
rect 423338 238294 453878 238350
rect 453934 238294 454002 238350
rect 454058 238294 484598 238350
rect 484654 238294 484722 238350
rect 484778 238294 515318 238350
rect 515374 238294 515442 238350
rect 515498 238294 546038 238350
rect 546094 238294 546162 238350
rect 546218 238294 561250 238350
rect 561306 238294 561374 238350
rect 561430 238294 561498 238350
rect 561554 238294 561622 238350
rect 561678 238294 579250 238350
rect 579306 238294 579374 238350
rect 579430 238294 579498 238350
rect 579554 238294 579622 238350
rect 579678 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597980 238350
rect -1916 238226 597980 238294
rect -1916 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 3250 238226
rect 3306 238170 3374 238226
rect 3430 238170 3498 238226
rect 3554 238170 3622 238226
rect 3678 238170 21250 238226
rect 21306 238170 21374 238226
rect 21430 238170 21498 238226
rect 21554 238170 21622 238226
rect 21678 238170 39250 238226
rect 39306 238170 39374 238226
rect 39430 238170 39498 238226
rect 39554 238170 39622 238226
rect 39678 238170 54518 238226
rect 54574 238170 54642 238226
rect 54698 238170 57250 238226
rect 57306 238170 57374 238226
rect 57430 238170 57498 238226
rect 57554 238170 57622 238226
rect 57678 238170 75250 238226
rect 75306 238170 75374 238226
rect 75430 238170 75498 238226
rect 75554 238170 75622 238226
rect 75678 238170 85238 238226
rect 85294 238170 85362 238226
rect 85418 238170 93250 238226
rect 93306 238170 93374 238226
rect 93430 238170 93498 238226
rect 93554 238170 93622 238226
rect 93678 238170 111250 238226
rect 111306 238170 111374 238226
rect 111430 238170 111498 238226
rect 111554 238170 111622 238226
rect 111678 238170 115958 238226
rect 116014 238170 116082 238226
rect 116138 238170 146678 238226
rect 146734 238170 146802 238226
rect 146858 238170 177398 238226
rect 177454 238170 177522 238226
rect 177578 238170 208118 238226
rect 208174 238170 208242 238226
rect 208298 238170 238838 238226
rect 238894 238170 238962 238226
rect 239018 238170 269558 238226
rect 269614 238170 269682 238226
rect 269738 238170 300278 238226
rect 300334 238170 300402 238226
rect 300458 238170 330998 238226
rect 331054 238170 331122 238226
rect 331178 238170 361718 238226
rect 361774 238170 361842 238226
rect 361898 238170 392438 238226
rect 392494 238170 392562 238226
rect 392618 238170 423158 238226
rect 423214 238170 423282 238226
rect 423338 238170 453878 238226
rect 453934 238170 454002 238226
rect 454058 238170 484598 238226
rect 484654 238170 484722 238226
rect 484778 238170 515318 238226
rect 515374 238170 515442 238226
rect 515498 238170 546038 238226
rect 546094 238170 546162 238226
rect 546218 238170 561250 238226
rect 561306 238170 561374 238226
rect 561430 238170 561498 238226
rect 561554 238170 561622 238226
rect 561678 238170 579250 238226
rect 579306 238170 579374 238226
rect 579430 238170 579498 238226
rect 579554 238170 579622 238226
rect 579678 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597980 238226
rect -1916 238102 597980 238170
rect -1916 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 3250 238102
rect 3306 238046 3374 238102
rect 3430 238046 3498 238102
rect 3554 238046 3622 238102
rect 3678 238046 21250 238102
rect 21306 238046 21374 238102
rect 21430 238046 21498 238102
rect 21554 238046 21622 238102
rect 21678 238046 39250 238102
rect 39306 238046 39374 238102
rect 39430 238046 39498 238102
rect 39554 238046 39622 238102
rect 39678 238046 54518 238102
rect 54574 238046 54642 238102
rect 54698 238046 57250 238102
rect 57306 238046 57374 238102
rect 57430 238046 57498 238102
rect 57554 238046 57622 238102
rect 57678 238046 75250 238102
rect 75306 238046 75374 238102
rect 75430 238046 75498 238102
rect 75554 238046 75622 238102
rect 75678 238046 85238 238102
rect 85294 238046 85362 238102
rect 85418 238046 93250 238102
rect 93306 238046 93374 238102
rect 93430 238046 93498 238102
rect 93554 238046 93622 238102
rect 93678 238046 111250 238102
rect 111306 238046 111374 238102
rect 111430 238046 111498 238102
rect 111554 238046 111622 238102
rect 111678 238046 115958 238102
rect 116014 238046 116082 238102
rect 116138 238046 146678 238102
rect 146734 238046 146802 238102
rect 146858 238046 177398 238102
rect 177454 238046 177522 238102
rect 177578 238046 208118 238102
rect 208174 238046 208242 238102
rect 208298 238046 238838 238102
rect 238894 238046 238962 238102
rect 239018 238046 269558 238102
rect 269614 238046 269682 238102
rect 269738 238046 300278 238102
rect 300334 238046 300402 238102
rect 300458 238046 330998 238102
rect 331054 238046 331122 238102
rect 331178 238046 361718 238102
rect 361774 238046 361842 238102
rect 361898 238046 392438 238102
rect 392494 238046 392562 238102
rect 392618 238046 423158 238102
rect 423214 238046 423282 238102
rect 423338 238046 453878 238102
rect 453934 238046 454002 238102
rect 454058 238046 484598 238102
rect 484654 238046 484722 238102
rect 484778 238046 515318 238102
rect 515374 238046 515442 238102
rect 515498 238046 546038 238102
rect 546094 238046 546162 238102
rect 546218 238046 561250 238102
rect 561306 238046 561374 238102
rect 561430 238046 561498 238102
rect 561554 238046 561622 238102
rect 561678 238046 579250 238102
rect 579306 238046 579374 238102
rect 579430 238046 579498 238102
rect 579554 238046 579622 238102
rect 579678 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597980 238102
rect -1916 237978 597980 238046
rect -1916 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 3250 237978
rect 3306 237922 3374 237978
rect 3430 237922 3498 237978
rect 3554 237922 3622 237978
rect 3678 237922 21250 237978
rect 21306 237922 21374 237978
rect 21430 237922 21498 237978
rect 21554 237922 21622 237978
rect 21678 237922 39250 237978
rect 39306 237922 39374 237978
rect 39430 237922 39498 237978
rect 39554 237922 39622 237978
rect 39678 237922 54518 237978
rect 54574 237922 54642 237978
rect 54698 237922 57250 237978
rect 57306 237922 57374 237978
rect 57430 237922 57498 237978
rect 57554 237922 57622 237978
rect 57678 237922 75250 237978
rect 75306 237922 75374 237978
rect 75430 237922 75498 237978
rect 75554 237922 75622 237978
rect 75678 237922 85238 237978
rect 85294 237922 85362 237978
rect 85418 237922 93250 237978
rect 93306 237922 93374 237978
rect 93430 237922 93498 237978
rect 93554 237922 93622 237978
rect 93678 237922 111250 237978
rect 111306 237922 111374 237978
rect 111430 237922 111498 237978
rect 111554 237922 111622 237978
rect 111678 237922 115958 237978
rect 116014 237922 116082 237978
rect 116138 237922 146678 237978
rect 146734 237922 146802 237978
rect 146858 237922 177398 237978
rect 177454 237922 177522 237978
rect 177578 237922 208118 237978
rect 208174 237922 208242 237978
rect 208298 237922 238838 237978
rect 238894 237922 238962 237978
rect 239018 237922 269558 237978
rect 269614 237922 269682 237978
rect 269738 237922 300278 237978
rect 300334 237922 300402 237978
rect 300458 237922 330998 237978
rect 331054 237922 331122 237978
rect 331178 237922 361718 237978
rect 361774 237922 361842 237978
rect 361898 237922 392438 237978
rect 392494 237922 392562 237978
rect 392618 237922 423158 237978
rect 423214 237922 423282 237978
rect 423338 237922 453878 237978
rect 453934 237922 454002 237978
rect 454058 237922 484598 237978
rect 484654 237922 484722 237978
rect 484778 237922 515318 237978
rect 515374 237922 515442 237978
rect 515498 237922 546038 237978
rect 546094 237922 546162 237978
rect 546218 237922 561250 237978
rect 561306 237922 561374 237978
rect 561430 237922 561498 237978
rect 561554 237922 561622 237978
rect 561678 237922 579250 237978
rect 579306 237922 579374 237978
rect 579430 237922 579498 237978
rect 579554 237922 579622 237978
rect 579678 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597980 237978
rect -1916 237826 597980 237922
rect -1916 226350 597980 226446
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 6970 226350
rect 7026 226294 7094 226350
rect 7150 226294 7218 226350
rect 7274 226294 7342 226350
rect 7398 226294 24970 226350
rect 25026 226294 25094 226350
rect 25150 226294 25218 226350
rect 25274 226294 25342 226350
rect 25398 226294 42970 226350
rect 43026 226294 43094 226350
rect 43150 226294 43218 226350
rect 43274 226294 43342 226350
rect 43398 226294 60970 226350
rect 61026 226294 61094 226350
rect 61150 226294 61218 226350
rect 61274 226294 61342 226350
rect 61398 226294 69878 226350
rect 69934 226294 70002 226350
rect 70058 226294 78970 226350
rect 79026 226294 79094 226350
rect 79150 226294 79218 226350
rect 79274 226294 79342 226350
rect 79398 226294 96970 226350
rect 97026 226294 97094 226350
rect 97150 226294 97218 226350
rect 97274 226294 97342 226350
rect 97398 226294 100598 226350
rect 100654 226294 100722 226350
rect 100778 226294 131318 226350
rect 131374 226294 131442 226350
rect 131498 226294 162038 226350
rect 162094 226294 162162 226350
rect 162218 226294 192758 226350
rect 192814 226294 192882 226350
rect 192938 226294 223478 226350
rect 223534 226294 223602 226350
rect 223658 226294 254198 226350
rect 254254 226294 254322 226350
rect 254378 226294 284918 226350
rect 284974 226294 285042 226350
rect 285098 226294 315638 226350
rect 315694 226294 315762 226350
rect 315818 226294 346358 226350
rect 346414 226294 346482 226350
rect 346538 226294 377078 226350
rect 377134 226294 377202 226350
rect 377258 226294 407798 226350
rect 407854 226294 407922 226350
rect 407978 226294 438518 226350
rect 438574 226294 438642 226350
rect 438698 226294 469238 226350
rect 469294 226294 469362 226350
rect 469418 226294 499958 226350
rect 500014 226294 500082 226350
rect 500138 226294 530678 226350
rect 530734 226294 530802 226350
rect 530858 226294 564970 226350
rect 565026 226294 565094 226350
rect 565150 226294 565218 226350
rect 565274 226294 565342 226350
rect 565398 226294 582970 226350
rect 583026 226294 583094 226350
rect 583150 226294 583218 226350
rect 583274 226294 583342 226350
rect 583398 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect -1916 226226 597980 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 6970 226226
rect 7026 226170 7094 226226
rect 7150 226170 7218 226226
rect 7274 226170 7342 226226
rect 7398 226170 24970 226226
rect 25026 226170 25094 226226
rect 25150 226170 25218 226226
rect 25274 226170 25342 226226
rect 25398 226170 42970 226226
rect 43026 226170 43094 226226
rect 43150 226170 43218 226226
rect 43274 226170 43342 226226
rect 43398 226170 60970 226226
rect 61026 226170 61094 226226
rect 61150 226170 61218 226226
rect 61274 226170 61342 226226
rect 61398 226170 69878 226226
rect 69934 226170 70002 226226
rect 70058 226170 78970 226226
rect 79026 226170 79094 226226
rect 79150 226170 79218 226226
rect 79274 226170 79342 226226
rect 79398 226170 96970 226226
rect 97026 226170 97094 226226
rect 97150 226170 97218 226226
rect 97274 226170 97342 226226
rect 97398 226170 100598 226226
rect 100654 226170 100722 226226
rect 100778 226170 131318 226226
rect 131374 226170 131442 226226
rect 131498 226170 162038 226226
rect 162094 226170 162162 226226
rect 162218 226170 192758 226226
rect 192814 226170 192882 226226
rect 192938 226170 223478 226226
rect 223534 226170 223602 226226
rect 223658 226170 254198 226226
rect 254254 226170 254322 226226
rect 254378 226170 284918 226226
rect 284974 226170 285042 226226
rect 285098 226170 315638 226226
rect 315694 226170 315762 226226
rect 315818 226170 346358 226226
rect 346414 226170 346482 226226
rect 346538 226170 377078 226226
rect 377134 226170 377202 226226
rect 377258 226170 407798 226226
rect 407854 226170 407922 226226
rect 407978 226170 438518 226226
rect 438574 226170 438642 226226
rect 438698 226170 469238 226226
rect 469294 226170 469362 226226
rect 469418 226170 499958 226226
rect 500014 226170 500082 226226
rect 500138 226170 530678 226226
rect 530734 226170 530802 226226
rect 530858 226170 564970 226226
rect 565026 226170 565094 226226
rect 565150 226170 565218 226226
rect 565274 226170 565342 226226
rect 565398 226170 582970 226226
rect 583026 226170 583094 226226
rect 583150 226170 583218 226226
rect 583274 226170 583342 226226
rect 583398 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect -1916 226102 597980 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 6970 226102
rect 7026 226046 7094 226102
rect 7150 226046 7218 226102
rect 7274 226046 7342 226102
rect 7398 226046 24970 226102
rect 25026 226046 25094 226102
rect 25150 226046 25218 226102
rect 25274 226046 25342 226102
rect 25398 226046 42970 226102
rect 43026 226046 43094 226102
rect 43150 226046 43218 226102
rect 43274 226046 43342 226102
rect 43398 226046 60970 226102
rect 61026 226046 61094 226102
rect 61150 226046 61218 226102
rect 61274 226046 61342 226102
rect 61398 226046 69878 226102
rect 69934 226046 70002 226102
rect 70058 226046 78970 226102
rect 79026 226046 79094 226102
rect 79150 226046 79218 226102
rect 79274 226046 79342 226102
rect 79398 226046 96970 226102
rect 97026 226046 97094 226102
rect 97150 226046 97218 226102
rect 97274 226046 97342 226102
rect 97398 226046 100598 226102
rect 100654 226046 100722 226102
rect 100778 226046 131318 226102
rect 131374 226046 131442 226102
rect 131498 226046 162038 226102
rect 162094 226046 162162 226102
rect 162218 226046 192758 226102
rect 192814 226046 192882 226102
rect 192938 226046 223478 226102
rect 223534 226046 223602 226102
rect 223658 226046 254198 226102
rect 254254 226046 254322 226102
rect 254378 226046 284918 226102
rect 284974 226046 285042 226102
rect 285098 226046 315638 226102
rect 315694 226046 315762 226102
rect 315818 226046 346358 226102
rect 346414 226046 346482 226102
rect 346538 226046 377078 226102
rect 377134 226046 377202 226102
rect 377258 226046 407798 226102
rect 407854 226046 407922 226102
rect 407978 226046 438518 226102
rect 438574 226046 438642 226102
rect 438698 226046 469238 226102
rect 469294 226046 469362 226102
rect 469418 226046 499958 226102
rect 500014 226046 500082 226102
rect 500138 226046 530678 226102
rect 530734 226046 530802 226102
rect 530858 226046 564970 226102
rect 565026 226046 565094 226102
rect 565150 226046 565218 226102
rect 565274 226046 565342 226102
rect 565398 226046 582970 226102
rect 583026 226046 583094 226102
rect 583150 226046 583218 226102
rect 583274 226046 583342 226102
rect 583398 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect -1916 225978 597980 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 6970 225978
rect 7026 225922 7094 225978
rect 7150 225922 7218 225978
rect 7274 225922 7342 225978
rect 7398 225922 24970 225978
rect 25026 225922 25094 225978
rect 25150 225922 25218 225978
rect 25274 225922 25342 225978
rect 25398 225922 42970 225978
rect 43026 225922 43094 225978
rect 43150 225922 43218 225978
rect 43274 225922 43342 225978
rect 43398 225922 60970 225978
rect 61026 225922 61094 225978
rect 61150 225922 61218 225978
rect 61274 225922 61342 225978
rect 61398 225922 69878 225978
rect 69934 225922 70002 225978
rect 70058 225922 78970 225978
rect 79026 225922 79094 225978
rect 79150 225922 79218 225978
rect 79274 225922 79342 225978
rect 79398 225922 96970 225978
rect 97026 225922 97094 225978
rect 97150 225922 97218 225978
rect 97274 225922 97342 225978
rect 97398 225922 100598 225978
rect 100654 225922 100722 225978
rect 100778 225922 131318 225978
rect 131374 225922 131442 225978
rect 131498 225922 162038 225978
rect 162094 225922 162162 225978
rect 162218 225922 192758 225978
rect 192814 225922 192882 225978
rect 192938 225922 223478 225978
rect 223534 225922 223602 225978
rect 223658 225922 254198 225978
rect 254254 225922 254322 225978
rect 254378 225922 284918 225978
rect 284974 225922 285042 225978
rect 285098 225922 315638 225978
rect 315694 225922 315762 225978
rect 315818 225922 346358 225978
rect 346414 225922 346482 225978
rect 346538 225922 377078 225978
rect 377134 225922 377202 225978
rect 377258 225922 407798 225978
rect 407854 225922 407922 225978
rect 407978 225922 438518 225978
rect 438574 225922 438642 225978
rect 438698 225922 469238 225978
rect 469294 225922 469362 225978
rect 469418 225922 499958 225978
rect 500014 225922 500082 225978
rect 500138 225922 530678 225978
rect 530734 225922 530802 225978
rect 530858 225922 564970 225978
rect 565026 225922 565094 225978
rect 565150 225922 565218 225978
rect 565274 225922 565342 225978
rect 565398 225922 582970 225978
rect 583026 225922 583094 225978
rect 583150 225922 583218 225978
rect 583274 225922 583342 225978
rect 583398 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect -1916 225826 597980 225922
rect -1916 220350 597980 220446
rect -1916 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 3250 220350
rect 3306 220294 3374 220350
rect 3430 220294 3498 220350
rect 3554 220294 3622 220350
rect 3678 220294 21250 220350
rect 21306 220294 21374 220350
rect 21430 220294 21498 220350
rect 21554 220294 21622 220350
rect 21678 220294 39250 220350
rect 39306 220294 39374 220350
rect 39430 220294 39498 220350
rect 39554 220294 39622 220350
rect 39678 220294 54518 220350
rect 54574 220294 54642 220350
rect 54698 220294 57250 220350
rect 57306 220294 57374 220350
rect 57430 220294 57498 220350
rect 57554 220294 57622 220350
rect 57678 220294 75250 220350
rect 75306 220294 75374 220350
rect 75430 220294 75498 220350
rect 75554 220294 75622 220350
rect 75678 220294 85238 220350
rect 85294 220294 85362 220350
rect 85418 220294 93250 220350
rect 93306 220294 93374 220350
rect 93430 220294 93498 220350
rect 93554 220294 93622 220350
rect 93678 220294 111250 220350
rect 111306 220294 111374 220350
rect 111430 220294 111498 220350
rect 111554 220294 111622 220350
rect 111678 220294 115958 220350
rect 116014 220294 116082 220350
rect 116138 220294 146678 220350
rect 146734 220294 146802 220350
rect 146858 220294 177398 220350
rect 177454 220294 177522 220350
rect 177578 220294 208118 220350
rect 208174 220294 208242 220350
rect 208298 220294 238838 220350
rect 238894 220294 238962 220350
rect 239018 220294 269558 220350
rect 269614 220294 269682 220350
rect 269738 220294 300278 220350
rect 300334 220294 300402 220350
rect 300458 220294 330998 220350
rect 331054 220294 331122 220350
rect 331178 220294 361718 220350
rect 361774 220294 361842 220350
rect 361898 220294 392438 220350
rect 392494 220294 392562 220350
rect 392618 220294 423158 220350
rect 423214 220294 423282 220350
rect 423338 220294 453878 220350
rect 453934 220294 454002 220350
rect 454058 220294 484598 220350
rect 484654 220294 484722 220350
rect 484778 220294 515318 220350
rect 515374 220294 515442 220350
rect 515498 220294 546038 220350
rect 546094 220294 546162 220350
rect 546218 220294 561250 220350
rect 561306 220294 561374 220350
rect 561430 220294 561498 220350
rect 561554 220294 561622 220350
rect 561678 220294 579250 220350
rect 579306 220294 579374 220350
rect 579430 220294 579498 220350
rect 579554 220294 579622 220350
rect 579678 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597980 220350
rect -1916 220226 597980 220294
rect -1916 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 3250 220226
rect 3306 220170 3374 220226
rect 3430 220170 3498 220226
rect 3554 220170 3622 220226
rect 3678 220170 21250 220226
rect 21306 220170 21374 220226
rect 21430 220170 21498 220226
rect 21554 220170 21622 220226
rect 21678 220170 39250 220226
rect 39306 220170 39374 220226
rect 39430 220170 39498 220226
rect 39554 220170 39622 220226
rect 39678 220170 54518 220226
rect 54574 220170 54642 220226
rect 54698 220170 57250 220226
rect 57306 220170 57374 220226
rect 57430 220170 57498 220226
rect 57554 220170 57622 220226
rect 57678 220170 75250 220226
rect 75306 220170 75374 220226
rect 75430 220170 75498 220226
rect 75554 220170 75622 220226
rect 75678 220170 85238 220226
rect 85294 220170 85362 220226
rect 85418 220170 93250 220226
rect 93306 220170 93374 220226
rect 93430 220170 93498 220226
rect 93554 220170 93622 220226
rect 93678 220170 111250 220226
rect 111306 220170 111374 220226
rect 111430 220170 111498 220226
rect 111554 220170 111622 220226
rect 111678 220170 115958 220226
rect 116014 220170 116082 220226
rect 116138 220170 146678 220226
rect 146734 220170 146802 220226
rect 146858 220170 177398 220226
rect 177454 220170 177522 220226
rect 177578 220170 208118 220226
rect 208174 220170 208242 220226
rect 208298 220170 238838 220226
rect 238894 220170 238962 220226
rect 239018 220170 269558 220226
rect 269614 220170 269682 220226
rect 269738 220170 300278 220226
rect 300334 220170 300402 220226
rect 300458 220170 330998 220226
rect 331054 220170 331122 220226
rect 331178 220170 361718 220226
rect 361774 220170 361842 220226
rect 361898 220170 392438 220226
rect 392494 220170 392562 220226
rect 392618 220170 423158 220226
rect 423214 220170 423282 220226
rect 423338 220170 453878 220226
rect 453934 220170 454002 220226
rect 454058 220170 484598 220226
rect 484654 220170 484722 220226
rect 484778 220170 515318 220226
rect 515374 220170 515442 220226
rect 515498 220170 546038 220226
rect 546094 220170 546162 220226
rect 546218 220170 561250 220226
rect 561306 220170 561374 220226
rect 561430 220170 561498 220226
rect 561554 220170 561622 220226
rect 561678 220170 579250 220226
rect 579306 220170 579374 220226
rect 579430 220170 579498 220226
rect 579554 220170 579622 220226
rect 579678 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597980 220226
rect -1916 220102 597980 220170
rect -1916 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 3250 220102
rect 3306 220046 3374 220102
rect 3430 220046 3498 220102
rect 3554 220046 3622 220102
rect 3678 220046 21250 220102
rect 21306 220046 21374 220102
rect 21430 220046 21498 220102
rect 21554 220046 21622 220102
rect 21678 220046 39250 220102
rect 39306 220046 39374 220102
rect 39430 220046 39498 220102
rect 39554 220046 39622 220102
rect 39678 220046 54518 220102
rect 54574 220046 54642 220102
rect 54698 220046 57250 220102
rect 57306 220046 57374 220102
rect 57430 220046 57498 220102
rect 57554 220046 57622 220102
rect 57678 220046 75250 220102
rect 75306 220046 75374 220102
rect 75430 220046 75498 220102
rect 75554 220046 75622 220102
rect 75678 220046 85238 220102
rect 85294 220046 85362 220102
rect 85418 220046 93250 220102
rect 93306 220046 93374 220102
rect 93430 220046 93498 220102
rect 93554 220046 93622 220102
rect 93678 220046 111250 220102
rect 111306 220046 111374 220102
rect 111430 220046 111498 220102
rect 111554 220046 111622 220102
rect 111678 220046 115958 220102
rect 116014 220046 116082 220102
rect 116138 220046 146678 220102
rect 146734 220046 146802 220102
rect 146858 220046 177398 220102
rect 177454 220046 177522 220102
rect 177578 220046 208118 220102
rect 208174 220046 208242 220102
rect 208298 220046 238838 220102
rect 238894 220046 238962 220102
rect 239018 220046 269558 220102
rect 269614 220046 269682 220102
rect 269738 220046 300278 220102
rect 300334 220046 300402 220102
rect 300458 220046 330998 220102
rect 331054 220046 331122 220102
rect 331178 220046 361718 220102
rect 361774 220046 361842 220102
rect 361898 220046 392438 220102
rect 392494 220046 392562 220102
rect 392618 220046 423158 220102
rect 423214 220046 423282 220102
rect 423338 220046 453878 220102
rect 453934 220046 454002 220102
rect 454058 220046 484598 220102
rect 484654 220046 484722 220102
rect 484778 220046 515318 220102
rect 515374 220046 515442 220102
rect 515498 220046 546038 220102
rect 546094 220046 546162 220102
rect 546218 220046 561250 220102
rect 561306 220046 561374 220102
rect 561430 220046 561498 220102
rect 561554 220046 561622 220102
rect 561678 220046 579250 220102
rect 579306 220046 579374 220102
rect 579430 220046 579498 220102
rect 579554 220046 579622 220102
rect 579678 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597980 220102
rect -1916 219978 597980 220046
rect -1916 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 3250 219978
rect 3306 219922 3374 219978
rect 3430 219922 3498 219978
rect 3554 219922 3622 219978
rect 3678 219922 21250 219978
rect 21306 219922 21374 219978
rect 21430 219922 21498 219978
rect 21554 219922 21622 219978
rect 21678 219922 39250 219978
rect 39306 219922 39374 219978
rect 39430 219922 39498 219978
rect 39554 219922 39622 219978
rect 39678 219922 54518 219978
rect 54574 219922 54642 219978
rect 54698 219922 57250 219978
rect 57306 219922 57374 219978
rect 57430 219922 57498 219978
rect 57554 219922 57622 219978
rect 57678 219922 75250 219978
rect 75306 219922 75374 219978
rect 75430 219922 75498 219978
rect 75554 219922 75622 219978
rect 75678 219922 85238 219978
rect 85294 219922 85362 219978
rect 85418 219922 93250 219978
rect 93306 219922 93374 219978
rect 93430 219922 93498 219978
rect 93554 219922 93622 219978
rect 93678 219922 111250 219978
rect 111306 219922 111374 219978
rect 111430 219922 111498 219978
rect 111554 219922 111622 219978
rect 111678 219922 115958 219978
rect 116014 219922 116082 219978
rect 116138 219922 146678 219978
rect 146734 219922 146802 219978
rect 146858 219922 177398 219978
rect 177454 219922 177522 219978
rect 177578 219922 208118 219978
rect 208174 219922 208242 219978
rect 208298 219922 238838 219978
rect 238894 219922 238962 219978
rect 239018 219922 269558 219978
rect 269614 219922 269682 219978
rect 269738 219922 300278 219978
rect 300334 219922 300402 219978
rect 300458 219922 330998 219978
rect 331054 219922 331122 219978
rect 331178 219922 361718 219978
rect 361774 219922 361842 219978
rect 361898 219922 392438 219978
rect 392494 219922 392562 219978
rect 392618 219922 423158 219978
rect 423214 219922 423282 219978
rect 423338 219922 453878 219978
rect 453934 219922 454002 219978
rect 454058 219922 484598 219978
rect 484654 219922 484722 219978
rect 484778 219922 515318 219978
rect 515374 219922 515442 219978
rect 515498 219922 546038 219978
rect 546094 219922 546162 219978
rect 546218 219922 561250 219978
rect 561306 219922 561374 219978
rect 561430 219922 561498 219978
rect 561554 219922 561622 219978
rect 561678 219922 579250 219978
rect 579306 219922 579374 219978
rect 579430 219922 579498 219978
rect 579554 219922 579622 219978
rect 579678 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597980 219978
rect -1916 219826 597980 219922
rect -1916 208350 597980 208446
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 6970 208350
rect 7026 208294 7094 208350
rect 7150 208294 7218 208350
rect 7274 208294 7342 208350
rect 7398 208294 24970 208350
rect 25026 208294 25094 208350
rect 25150 208294 25218 208350
rect 25274 208294 25342 208350
rect 25398 208294 42970 208350
rect 43026 208294 43094 208350
rect 43150 208294 43218 208350
rect 43274 208294 43342 208350
rect 43398 208294 60970 208350
rect 61026 208294 61094 208350
rect 61150 208294 61218 208350
rect 61274 208294 61342 208350
rect 61398 208294 69878 208350
rect 69934 208294 70002 208350
rect 70058 208294 78970 208350
rect 79026 208294 79094 208350
rect 79150 208294 79218 208350
rect 79274 208294 79342 208350
rect 79398 208294 96970 208350
rect 97026 208294 97094 208350
rect 97150 208294 97218 208350
rect 97274 208294 97342 208350
rect 97398 208294 100598 208350
rect 100654 208294 100722 208350
rect 100778 208294 131318 208350
rect 131374 208294 131442 208350
rect 131498 208294 162038 208350
rect 162094 208294 162162 208350
rect 162218 208294 192758 208350
rect 192814 208294 192882 208350
rect 192938 208294 223478 208350
rect 223534 208294 223602 208350
rect 223658 208294 254198 208350
rect 254254 208294 254322 208350
rect 254378 208294 284918 208350
rect 284974 208294 285042 208350
rect 285098 208294 315638 208350
rect 315694 208294 315762 208350
rect 315818 208294 346358 208350
rect 346414 208294 346482 208350
rect 346538 208294 377078 208350
rect 377134 208294 377202 208350
rect 377258 208294 407798 208350
rect 407854 208294 407922 208350
rect 407978 208294 438518 208350
rect 438574 208294 438642 208350
rect 438698 208294 469238 208350
rect 469294 208294 469362 208350
rect 469418 208294 499958 208350
rect 500014 208294 500082 208350
rect 500138 208294 530678 208350
rect 530734 208294 530802 208350
rect 530858 208294 564970 208350
rect 565026 208294 565094 208350
rect 565150 208294 565218 208350
rect 565274 208294 565342 208350
rect 565398 208294 582970 208350
rect 583026 208294 583094 208350
rect 583150 208294 583218 208350
rect 583274 208294 583342 208350
rect 583398 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect -1916 208226 597980 208294
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 6970 208226
rect 7026 208170 7094 208226
rect 7150 208170 7218 208226
rect 7274 208170 7342 208226
rect 7398 208170 24970 208226
rect 25026 208170 25094 208226
rect 25150 208170 25218 208226
rect 25274 208170 25342 208226
rect 25398 208170 42970 208226
rect 43026 208170 43094 208226
rect 43150 208170 43218 208226
rect 43274 208170 43342 208226
rect 43398 208170 60970 208226
rect 61026 208170 61094 208226
rect 61150 208170 61218 208226
rect 61274 208170 61342 208226
rect 61398 208170 69878 208226
rect 69934 208170 70002 208226
rect 70058 208170 78970 208226
rect 79026 208170 79094 208226
rect 79150 208170 79218 208226
rect 79274 208170 79342 208226
rect 79398 208170 96970 208226
rect 97026 208170 97094 208226
rect 97150 208170 97218 208226
rect 97274 208170 97342 208226
rect 97398 208170 100598 208226
rect 100654 208170 100722 208226
rect 100778 208170 131318 208226
rect 131374 208170 131442 208226
rect 131498 208170 162038 208226
rect 162094 208170 162162 208226
rect 162218 208170 192758 208226
rect 192814 208170 192882 208226
rect 192938 208170 223478 208226
rect 223534 208170 223602 208226
rect 223658 208170 254198 208226
rect 254254 208170 254322 208226
rect 254378 208170 284918 208226
rect 284974 208170 285042 208226
rect 285098 208170 315638 208226
rect 315694 208170 315762 208226
rect 315818 208170 346358 208226
rect 346414 208170 346482 208226
rect 346538 208170 377078 208226
rect 377134 208170 377202 208226
rect 377258 208170 407798 208226
rect 407854 208170 407922 208226
rect 407978 208170 438518 208226
rect 438574 208170 438642 208226
rect 438698 208170 469238 208226
rect 469294 208170 469362 208226
rect 469418 208170 499958 208226
rect 500014 208170 500082 208226
rect 500138 208170 530678 208226
rect 530734 208170 530802 208226
rect 530858 208170 564970 208226
rect 565026 208170 565094 208226
rect 565150 208170 565218 208226
rect 565274 208170 565342 208226
rect 565398 208170 582970 208226
rect 583026 208170 583094 208226
rect 583150 208170 583218 208226
rect 583274 208170 583342 208226
rect 583398 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect -1916 208102 597980 208170
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 6970 208102
rect 7026 208046 7094 208102
rect 7150 208046 7218 208102
rect 7274 208046 7342 208102
rect 7398 208046 24970 208102
rect 25026 208046 25094 208102
rect 25150 208046 25218 208102
rect 25274 208046 25342 208102
rect 25398 208046 42970 208102
rect 43026 208046 43094 208102
rect 43150 208046 43218 208102
rect 43274 208046 43342 208102
rect 43398 208046 60970 208102
rect 61026 208046 61094 208102
rect 61150 208046 61218 208102
rect 61274 208046 61342 208102
rect 61398 208046 69878 208102
rect 69934 208046 70002 208102
rect 70058 208046 78970 208102
rect 79026 208046 79094 208102
rect 79150 208046 79218 208102
rect 79274 208046 79342 208102
rect 79398 208046 96970 208102
rect 97026 208046 97094 208102
rect 97150 208046 97218 208102
rect 97274 208046 97342 208102
rect 97398 208046 100598 208102
rect 100654 208046 100722 208102
rect 100778 208046 131318 208102
rect 131374 208046 131442 208102
rect 131498 208046 162038 208102
rect 162094 208046 162162 208102
rect 162218 208046 192758 208102
rect 192814 208046 192882 208102
rect 192938 208046 223478 208102
rect 223534 208046 223602 208102
rect 223658 208046 254198 208102
rect 254254 208046 254322 208102
rect 254378 208046 284918 208102
rect 284974 208046 285042 208102
rect 285098 208046 315638 208102
rect 315694 208046 315762 208102
rect 315818 208046 346358 208102
rect 346414 208046 346482 208102
rect 346538 208046 377078 208102
rect 377134 208046 377202 208102
rect 377258 208046 407798 208102
rect 407854 208046 407922 208102
rect 407978 208046 438518 208102
rect 438574 208046 438642 208102
rect 438698 208046 469238 208102
rect 469294 208046 469362 208102
rect 469418 208046 499958 208102
rect 500014 208046 500082 208102
rect 500138 208046 530678 208102
rect 530734 208046 530802 208102
rect 530858 208046 564970 208102
rect 565026 208046 565094 208102
rect 565150 208046 565218 208102
rect 565274 208046 565342 208102
rect 565398 208046 582970 208102
rect 583026 208046 583094 208102
rect 583150 208046 583218 208102
rect 583274 208046 583342 208102
rect 583398 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect -1916 207978 597980 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 6970 207978
rect 7026 207922 7094 207978
rect 7150 207922 7218 207978
rect 7274 207922 7342 207978
rect 7398 207922 24970 207978
rect 25026 207922 25094 207978
rect 25150 207922 25218 207978
rect 25274 207922 25342 207978
rect 25398 207922 42970 207978
rect 43026 207922 43094 207978
rect 43150 207922 43218 207978
rect 43274 207922 43342 207978
rect 43398 207922 60970 207978
rect 61026 207922 61094 207978
rect 61150 207922 61218 207978
rect 61274 207922 61342 207978
rect 61398 207922 69878 207978
rect 69934 207922 70002 207978
rect 70058 207922 78970 207978
rect 79026 207922 79094 207978
rect 79150 207922 79218 207978
rect 79274 207922 79342 207978
rect 79398 207922 96970 207978
rect 97026 207922 97094 207978
rect 97150 207922 97218 207978
rect 97274 207922 97342 207978
rect 97398 207922 100598 207978
rect 100654 207922 100722 207978
rect 100778 207922 131318 207978
rect 131374 207922 131442 207978
rect 131498 207922 162038 207978
rect 162094 207922 162162 207978
rect 162218 207922 192758 207978
rect 192814 207922 192882 207978
rect 192938 207922 223478 207978
rect 223534 207922 223602 207978
rect 223658 207922 254198 207978
rect 254254 207922 254322 207978
rect 254378 207922 284918 207978
rect 284974 207922 285042 207978
rect 285098 207922 315638 207978
rect 315694 207922 315762 207978
rect 315818 207922 346358 207978
rect 346414 207922 346482 207978
rect 346538 207922 377078 207978
rect 377134 207922 377202 207978
rect 377258 207922 407798 207978
rect 407854 207922 407922 207978
rect 407978 207922 438518 207978
rect 438574 207922 438642 207978
rect 438698 207922 469238 207978
rect 469294 207922 469362 207978
rect 469418 207922 499958 207978
rect 500014 207922 500082 207978
rect 500138 207922 530678 207978
rect 530734 207922 530802 207978
rect 530858 207922 564970 207978
rect 565026 207922 565094 207978
rect 565150 207922 565218 207978
rect 565274 207922 565342 207978
rect 565398 207922 582970 207978
rect 583026 207922 583094 207978
rect 583150 207922 583218 207978
rect 583274 207922 583342 207978
rect 583398 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect -1916 207826 597980 207922
rect -1916 202350 597980 202446
rect -1916 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 3250 202350
rect 3306 202294 3374 202350
rect 3430 202294 3498 202350
rect 3554 202294 3622 202350
rect 3678 202294 21250 202350
rect 21306 202294 21374 202350
rect 21430 202294 21498 202350
rect 21554 202294 21622 202350
rect 21678 202294 39250 202350
rect 39306 202294 39374 202350
rect 39430 202294 39498 202350
rect 39554 202294 39622 202350
rect 39678 202294 54518 202350
rect 54574 202294 54642 202350
rect 54698 202294 57250 202350
rect 57306 202294 57374 202350
rect 57430 202294 57498 202350
rect 57554 202294 57622 202350
rect 57678 202294 75250 202350
rect 75306 202294 75374 202350
rect 75430 202294 75498 202350
rect 75554 202294 75622 202350
rect 75678 202294 85238 202350
rect 85294 202294 85362 202350
rect 85418 202294 93250 202350
rect 93306 202294 93374 202350
rect 93430 202294 93498 202350
rect 93554 202294 93622 202350
rect 93678 202294 111250 202350
rect 111306 202294 111374 202350
rect 111430 202294 111498 202350
rect 111554 202294 111622 202350
rect 111678 202294 115958 202350
rect 116014 202294 116082 202350
rect 116138 202294 146678 202350
rect 146734 202294 146802 202350
rect 146858 202294 177398 202350
rect 177454 202294 177522 202350
rect 177578 202294 208118 202350
rect 208174 202294 208242 202350
rect 208298 202294 238838 202350
rect 238894 202294 238962 202350
rect 239018 202294 269558 202350
rect 269614 202294 269682 202350
rect 269738 202294 300278 202350
rect 300334 202294 300402 202350
rect 300458 202294 330998 202350
rect 331054 202294 331122 202350
rect 331178 202294 361718 202350
rect 361774 202294 361842 202350
rect 361898 202294 392438 202350
rect 392494 202294 392562 202350
rect 392618 202294 423158 202350
rect 423214 202294 423282 202350
rect 423338 202294 453878 202350
rect 453934 202294 454002 202350
rect 454058 202294 484598 202350
rect 484654 202294 484722 202350
rect 484778 202294 515318 202350
rect 515374 202294 515442 202350
rect 515498 202294 546038 202350
rect 546094 202294 546162 202350
rect 546218 202294 561250 202350
rect 561306 202294 561374 202350
rect 561430 202294 561498 202350
rect 561554 202294 561622 202350
rect 561678 202294 579250 202350
rect 579306 202294 579374 202350
rect 579430 202294 579498 202350
rect 579554 202294 579622 202350
rect 579678 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597980 202350
rect -1916 202226 597980 202294
rect -1916 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 3250 202226
rect 3306 202170 3374 202226
rect 3430 202170 3498 202226
rect 3554 202170 3622 202226
rect 3678 202170 21250 202226
rect 21306 202170 21374 202226
rect 21430 202170 21498 202226
rect 21554 202170 21622 202226
rect 21678 202170 39250 202226
rect 39306 202170 39374 202226
rect 39430 202170 39498 202226
rect 39554 202170 39622 202226
rect 39678 202170 54518 202226
rect 54574 202170 54642 202226
rect 54698 202170 57250 202226
rect 57306 202170 57374 202226
rect 57430 202170 57498 202226
rect 57554 202170 57622 202226
rect 57678 202170 75250 202226
rect 75306 202170 75374 202226
rect 75430 202170 75498 202226
rect 75554 202170 75622 202226
rect 75678 202170 85238 202226
rect 85294 202170 85362 202226
rect 85418 202170 93250 202226
rect 93306 202170 93374 202226
rect 93430 202170 93498 202226
rect 93554 202170 93622 202226
rect 93678 202170 111250 202226
rect 111306 202170 111374 202226
rect 111430 202170 111498 202226
rect 111554 202170 111622 202226
rect 111678 202170 115958 202226
rect 116014 202170 116082 202226
rect 116138 202170 146678 202226
rect 146734 202170 146802 202226
rect 146858 202170 177398 202226
rect 177454 202170 177522 202226
rect 177578 202170 208118 202226
rect 208174 202170 208242 202226
rect 208298 202170 238838 202226
rect 238894 202170 238962 202226
rect 239018 202170 269558 202226
rect 269614 202170 269682 202226
rect 269738 202170 300278 202226
rect 300334 202170 300402 202226
rect 300458 202170 330998 202226
rect 331054 202170 331122 202226
rect 331178 202170 361718 202226
rect 361774 202170 361842 202226
rect 361898 202170 392438 202226
rect 392494 202170 392562 202226
rect 392618 202170 423158 202226
rect 423214 202170 423282 202226
rect 423338 202170 453878 202226
rect 453934 202170 454002 202226
rect 454058 202170 484598 202226
rect 484654 202170 484722 202226
rect 484778 202170 515318 202226
rect 515374 202170 515442 202226
rect 515498 202170 546038 202226
rect 546094 202170 546162 202226
rect 546218 202170 561250 202226
rect 561306 202170 561374 202226
rect 561430 202170 561498 202226
rect 561554 202170 561622 202226
rect 561678 202170 579250 202226
rect 579306 202170 579374 202226
rect 579430 202170 579498 202226
rect 579554 202170 579622 202226
rect 579678 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597980 202226
rect -1916 202102 597980 202170
rect -1916 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 3250 202102
rect 3306 202046 3374 202102
rect 3430 202046 3498 202102
rect 3554 202046 3622 202102
rect 3678 202046 21250 202102
rect 21306 202046 21374 202102
rect 21430 202046 21498 202102
rect 21554 202046 21622 202102
rect 21678 202046 39250 202102
rect 39306 202046 39374 202102
rect 39430 202046 39498 202102
rect 39554 202046 39622 202102
rect 39678 202046 54518 202102
rect 54574 202046 54642 202102
rect 54698 202046 57250 202102
rect 57306 202046 57374 202102
rect 57430 202046 57498 202102
rect 57554 202046 57622 202102
rect 57678 202046 75250 202102
rect 75306 202046 75374 202102
rect 75430 202046 75498 202102
rect 75554 202046 75622 202102
rect 75678 202046 85238 202102
rect 85294 202046 85362 202102
rect 85418 202046 93250 202102
rect 93306 202046 93374 202102
rect 93430 202046 93498 202102
rect 93554 202046 93622 202102
rect 93678 202046 111250 202102
rect 111306 202046 111374 202102
rect 111430 202046 111498 202102
rect 111554 202046 111622 202102
rect 111678 202046 115958 202102
rect 116014 202046 116082 202102
rect 116138 202046 146678 202102
rect 146734 202046 146802 202102
rect 146858 202046 177398 202102
rect 177454 202046 177522 202102
rect 177578 202046 208118 202102
rect 208174 202046 208242 202102
rect 208298 202046 238838 202102
rect 238894 202046 238962 202102
rect 239018 202046 269558 202102
rect 269614 202046 269682 202102
rect 269738 202046 300278 202102
rect 300334 202046 300402 202102
rect 300458 202046 330998 202102
rect 331054 202046 331122 202102
rect 331178 202046 361718 202102
rect 361774 202046 361842 202102
rect 361898 202046 392438 202102
rect 392494 202046 392562 202102
rect 392618 202046 423158 202102
rect 423214 202046 423282 202102
rect 423338 202046 453878 202102
rect 453934 202046 454002 202102
rect 454058 202046 484598 202102
rect 484654 202046 484722 202102
rect 484778 202046 515318 202102
rect 515374 202046 515442 202102
rect 515498 202046 546038 202102
rect 546094 202046 546162 202102
rect 546218 202046 561250 202102
rect 561306 202046 561374 202102
rect 561430 202046 561498 202102
rect 561554 202046 561622 202102
rect 561678 202046 579250 202102
rect 579306 202046 579374 202102
rect 579430 202046 579498 202102
rect 579554 202046 579622 202102
rect 579678 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597980 202102
rect -1916 201978 597980 202046
rect -1916 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 3250 201978
rect 3306 201922 3374 201978
rect 3430 201922 3498 201978
rect 3554 201922 3622 201978
rect 3678 201922 21250 201978
rect 21306 201922 21374 201978
rect 21430 201922 21498 201978
rect 21554 201922 21622 201978
rect 21678 201922 39250 201978
rect 39306 201922 39374 201978
rect 39430 201922 39498 201978
rect 39554 201922 39622 201978
rect 39678 201922 54518 201978
rect 54574 201922 54642 201978
rect 54698 201922 57250 201978
rect 57306 201922 57374 201978
rect 57430 201922 57498 201978
rect 57554 201922 57622 201978
rect 57678 201922 75250 201978
rect 75306 201922 75374 201978
rect 75430 201922 75498 201978
rect 75554 201922 75622 201978
rect 75678 201922 85238 201978
rect 85294 201922 85362 201978
rect 85418 201922 93250 201978
rect 93306 201922 93374 201978
rect 93430 201922 93498 201978
rect 93554 201922 93622 201978
rect 93678 201922 111250 201978
rect 111306 201922 111374 201978
rect 111430 201922 111498 201978
rect 111554 201922 111622 201978
rect 111678 201922 115958 201978
rect 116014 201922 116082 201978
rect 116138 201922 146678 201978
rect 146734 201922 146802 201978
rect 146858 201922 177398 201978
rect 177454 201922 177522 201978
rect 177578 201922 208118 201978
rect 208174 201922 208242 201978
rect 208298 201922 238838 201978
rect 238894 201922 238962 201978
rect 239018 201922 269558 201978
rect 269614 201922 269682 201978
rect 269738 201922 300278 201978
rect 300334 201922 300402 201978
rect 300458 201922 330998 201978
rect 331054 201922 331122 201978
rect 331178 201922 361718 201978
rect 361774 201922 361842 201978
rect 361898 201922 392438 201978
rect 392494 201922 392562 201978
rect 392618 201922 423158 201978
rect 423214 201922 423282 201978
rect 423338 201922 453878 201978
rect 453934 201922 454002 201978
rect 454058 201922 484598 201978
rect 484654 201922 484722 201978
rect 484778 201922 515318 201978
rect 515374 201922 515442 201978
rect 515498 201922 546038 201978
rect 546094 201922 546162 201978
rect 546218 201922 561250 201978
rect 561306 201922 561374 201978
rect 561430 201922 561498 201978
rect 561554 201922 561622 201978
rect 561678 201922 579250 201978
rect 579306 201922 579374 201978
rect 579430 201922 579498 201978
rect 579554 201922 579622 201978
rect 579678 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597980 201978
rect -1916 201826 597980 201922
rect -1916 190350 597980 190446
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 6970 190350
rect 7026 190294 7094 190350
rect 7150 190294 7218 190350
rect 7274 190294 7342 190350
rect 7398 190294 24970 190350
rect 25026 190294 25094 190350
rect 25150 190294 25218 190350
rect 25274 190294 25342 190350
rect 25398 190294 42970 190350
rect 43026 190294 43094 190350
rect 43150 190294 43218 190350
rect 43274 190294 43342 190350
rect 43398 190294 60970 190350
rect 61026 190294 61094 190350
rect 61150 190294 61218 190350
rect 61274 190294 61342 190350
rect 61398 190294 69878 190350
rect 69934 190294 70002 190350
rect 70058 190294 78970 190350
rect 79026 190294 79094 190350
rect 79150 190294 79218 190350
rect 79274 190294 79342 190350
rect 79398 190294 96970 190350
rect 97026 190294 97094 190350
rect 97150 190294 97218 190350
rect 97274 190294 97342 190350
rect 97398 190294 100598 190350
rect 100654 190294 100722 190350
rect 100778 190294 131318 190350
rect 131374 190294 131442 190350
rect 131498 190294 162038 190350
rect 162094 190294 162162 190350
rect 162218 190294 192758 190350
rect 192814 190294 192882 190350
rect 192938 190294 223478 190350
rect 223534 190294 223602 190350
rect 223658 190294 254198 190350
rect 254254 190294 254322 190350
rect 254378 190294 284918 190350
rect 284974 190294 285042 190350
rect 285098 190294 315638 190350
rect 315694 190294 315762 190350
rect 315818 190294 346358 190350
rect 346414 190294 346482 190350
rect 346538 190294 377078 190350
rect 377134 190294 377202 190350
rect 377258 190294 407798 190350
rect 407854 190294 407922 190350
rect 407978 190294 438518 190350
rect 438574 190294 438642 190350
rect 438698 190294 469238 190350
rect 469294 190294 469362 190350
rect 469418 190294 499958 190350
rect 500014 190294 500082 190350
rect 500138 190294 530678 190350
rect 530734 190294 530802 190350
rect 530858 190294 564970 190350
rect 565026 190294 565094 190350
rect 565150 190294 565218 190350
rect 565274 190294 565342 190350
rect 565398 190294 582970 190350
rect 583026 190294 583094 190350
rect 583150 190294 583218 190350
rect 583274 190294 583342 190350
rect 583398 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect -1916 190226 597980 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 6970 190226
rect 7026 190170 7094 190226
rect 7150 190170 7218 190226
rect 7274 190170 7342 190226
rect 7398 190170 24970 190226
rect 25026 190170 25094 190226
rect 25150 190170 25218 190226
rect 25274 190170 25342 190226
rect 25398 190170 42970 190226
rect 43026 190170 43094 190226
rect 43150 190170 43218 190226
rect 43274 190170 43342 190226
rect 43398 190170 60970 190226
rect 61026 190170 61094 190226
rect 61150 190170 61218 190226
rect 61274 190170 61342 190226
rect 61398 190170 69878 190226
rect 69934 190170 70002 190226
rect 70058 190170 78970 190226
rect 79026 190170 79094 190226
rect 79150 190170 79218 190226
rect 79274 190170 79342 190226
rect 79398 190170 96970 190226
rect 97026 190170 97094 190226
rect 97150 190170 97218 190226
rect 97274 190170 97342 190226
rect 97398 190170 100598 190226
rect 100654 190170 100722 190226
rect 100778 190170 131318 190226
rect 131374 190170 131442 190226
rect 131498 190170 162038 190226
rect 162094 190170 162162 190226
rect 162218 190170 192758 190226
rect 192814 190170 192882 190226
rect 192938 190170 223478 190226
rect 223534 190170 223602 190226
rect 223658 190170 254198 190226
rect 254254 190170 254322 190226
rect 254378 190170 284918 190226
rect 284974 190170 285042 190226
rect 285098 190170 315638 190226
rect 315694 190170 315762 190226
rect 315818 190170 346358 190226
rect 346414 190170 346482 190226
rect 346538 190170 377078 190226
rect 377134 190170 377202 190226
rect 377258 190170 407798 190226
rect 407854 190170 407922 190226
rect 407978 190170 438518 190226
rect 438574 190170 438642 190226
rect 438698 190170 469238 190226
rect 469294 190170 469362 190226
rect 469418 190170 499958 190226
rect 500014 190170 500082 190226
rect 500138 190170 530678 190226
rect 530734 190170 530802 190226
rect 530858 190170 564970 190226
rect 565026 190170 565094 190226
rect 565150 190170 565218 190226
rect 565274 190170 565342 190226
rect 565398 190170 582970 190226
rect 583026 190170 583094 190226
rect 583150 190170 583218 190226
rect 583274 190170 583342 190226
rect 583398 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect -1916 190102 597980 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 6970 190102
rect 7026 190046 7094 190102
rect 7150 190046 7218 190102
rect 7274 190046 7342 190102
rect 7398 190046 24970 190102
rect 25026 190046 25094 190102
rect 25150 190046 25218 190102
rect 25274 190046 25342 190102
rect 25398 190046 42970 190102
rect 43026 190046 43094 190102
rect 43150 190046 43218 190102
rect 43274 190046 43342 190102
rect 43398 190046 60970 190102
rect 61026 190046 61094 190102
rect 61150 190046 61218 190102
rect 61274 190046 61342 190102
rect 61398 190046 69878 190102
rect 69934 190046 70002 190102
rect 70058 190046 78970 190102
rect 79026 190046 79094 190102
rect 79150 190046 79218 190102
rect 79274 190046 79342 190102
rect 79398 190046 96970 190102
rect 97026 190046 97094 190102
rect 97150 190046 97218 190102
rect 97274 190046 97342 190102
rect 97398 190046 100598 190102
rect 100654 190046 100722 190102
rect 100778 190046 131318 190102
rect 131374 190046 131442 190102
rect 131498 190046 162038 190102
rect 162094 190046 162162 190102
rect 162218 190046 192758 190102
rect 192814 190046 192882 190102
rect 192938 190046 223478 190102
rect 223534 190046 223602 190102
rect 223658 190046 254198 190102
rect 254254 190046 254322 190102
rect 254378 190046 284918 190102
rect 284974 190046 285042 190102
rect 285098 190046 315638 190102
rect 315694 190046 315762 190102
rect 315818 190046 346358 190102
rect 346414 190046 346482 190102
rect 346538 190046 377078 190102
rect 377134 190046 377202 190102
rect 377258 190046 407798 190102
rect 407854 190046 407922 190102
rect 407978 190046 438518 190102
rect 438574 190046 438642 190102
rect 438698 190046 469238 190102
rect 469294 190046 469362 190102
rect 469418 190046 499958 190102
rect 500014 190046 500082 190102
rect 500138 190046 530678 190102
rect 530734 190046 530802 190102
rect 530858 190046 564970 190102
rect 565026 190046 565094 190102
rect 565150 190046 565218 190102
rect 565274 190046 565342 190102
rect 565398 190046 582970 190102
rect 583026 190046 583094 190102
rect 583150 190046 583218 190102
rect 583274 190046 583342 190102
rect 583398 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect -1916 189978 597980 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 6970 189978
rect 7026 189922 7094 189978
rect 7150 189922 7218 189978
rect 7274 189922 7342 189978
rect 7398 189922 24970 189978
rect 25026 189922 25094 189978
rect 25150 189922 25218 189978
rect 25274 189922 25342 189978
rect 25398 189922 42970 189978
rect 43026 189922 43094 189978
rect 43150 189922 43218 189978
rect 43274 189922 43342 189978
rect 43398 189922 60970 189978
rect 61026 189922 61094 189978
rect 61150 189922 61218 189978
rect 61274 189922 61342 189978
rect 61398 189922 69878 189978
rect 69934 189922 70002 189978
rect 70058 189922 78970 189978
rect 79026 189922 79094 189978
rect 79150 189922 79218 189978
rect 79274 189922 79342 189978
rect 79398 189922 96970 189978
rect 97026 189922 97094 189978
rect 97150 189922 97218 189978
rect 97274 189922 97342 189978
rect 97398 189922 100598 189978
rect 100654 189922 100722 189978
rect 100778 189922 131318 189978
rect 131374 189922 131442 189978
rect 131498 189922 162038 189978
rect 162094 189922 162162 189978
rect 162218 189922 192758 189978
rect 192814 189922 192882 189978
rect 192938 189922 223478 189978
rect 223534 189922 223602 189978
rect 223658 189922 254198 189978
rect 254254 189922 254322 189978
rect 254378 189922 284918 189978
rect 284974 189922 285042 189978
rect 285098 189922 315638 189978
rect 315694 189922 315762 189978
rect 315818 189922 346358 189978
rect 346414 189922 346482 189978
rect 346538 189922 377078 189978
rect 377134 189922 377202 189978
rect 377258 189922 407798 189978
rect 407854 189922 407922 189978
rect 407978 189922 438518 189978
rect 438574 189922 438642 189978
rect 438698 189922 469238 189978
rect 469294 189922 469362 189978
rect 469418 189922 499958 189978
rect 500014 189922 500082 189978
rect 500138 189922 530678 189978
rect 530734 189922 530802 189978
rect 530858 189922 564970 189978
rect 565026 189922 565094 189978
rect 565150 189922 565218 189978
rect 565274 189922 565342 189978
rect 565398 189922 582970 189978
rect 583026 189922 583094 189978
rect 583150 189922 583218 189978
rect 583274 189922 583342 189978
rect 583398 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect -1916 189826 597980 189922
rect -1916 184350 597980 184446
rect -1916 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 3250 184350
rect 3306 184294 3374 184350
rect 3430 184294 3498 184350
rect 3554 184294 3622 184350
rect 3678 184294 21250 184350
rect 21306 184294 21374 184350
rect 21430 184294 21498 184350
rect 21554 184294 21622 184350
rect 21678 184294 39250 184350
rect 39306 184294 39374 184350
rect 39430 184294 39498 184350
rect 39554 184294 39622 184350
rect 39678 184294 54518 184350
rect 54574 184294 54642 184350
rect 54698 184294 57250 184350
rect 57306 184294 57374 184350
rect 57430 184294 57498 184350
rect 57554 184294 57622 184350
rect 57678 184294 75250 184350
rect 75306 184294 75374 184350
rect 75430 184294 75498 184350
rect 75554 184294 75622 184350
rect 75678 184294 85238 184350
rect 85294 184294 85362 184350
rect 85418 184294 93250 184350
rect 93306 184294 93374 184350
rect 93430 184294 93498 184350
rect 93554 184294 93622 184350
rect 93678 184294 111250 184350
rect 111306 184294 111374 184350
rect 111430 184294 111498 184350
rect 111554 184294 111622 184350
rect 111678 184294 115958 184350
rect 116014 184294 116082 184350
rect 116138 184294 146678 184350
rect 146734 184294 146802 184350
rect 146858 184294 177398 184350
rect 177454 184294 177522 184350
rect 177578 184294 208118 184350
rect 208174 184294 208242 184350
rect 208298 184294 238838 184350
rect 238894 184294 238962 184350
rect 239018 184294 269558 184350
rect 269614 184294 269682 184350
rect 269738 184294 300278 184350
rect 300334 184294 300402 184350
rect 300458 184294 330998 184350
rect 331054 184294 331122 184350
rect 331178 184294 361718 184350
rect 361774 184294 361842 184350
rect 361898 184294 392438 184350
rect 392494 184294 392562 184350
rect 392618 184294 423158 184350
rect 423214 184294 423282 184350
rect 423338 184294 453878 184350
rect 453934 184294 454002 184350
rect 454058 184294 484598 184350
rect 484654 184294 484722 184350
rect 484778 184294 515318 184350
rect 515374 184294 515442 184350
rect 515498 184294 546038 184350
rect 546094 184294 546162 184350
rect 546218 184294 561250 184350
rect 561306 184294 561374 184350
rect 561430 184294 561498 184350
rect 561554 184294 561622 184350
rect 561678 184294 579250 184350
rect 579306 184294 579374 184350
rect 579430 184294 579498 184350
rect 579554 184294 579622 184350
rect 579678 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597980 184350
rect -1916 184226 597980 184294
rect -1916 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 3250 184226
rect 3306 184170 3374 184226
rect 3430 184170 3498 184226
rect 3554 184170 3622 184226
rect 3678 184170 21250 184226
rect 21306 184170 21374 184226
rect 21430 184170 21498 184226
rect 21554 184170 21622 184226
rect 21678 184170 39250 184226
rect 39306 184170 39374 184226
rect 39430 184170 39498 184226
rect 39554 184170 39622 184226
rect 39678 184170 54518 184226
rect 54574 184170 54642 184226
rect 54698 184170 57250 184226
rect 57306 184170 57374 184226
rect 57430 184170 57498 184226
rect 57554 184170 57622 184226
rect 57678 184170 75250 184226
rect 75306 184170 75374 184226
rect 75430 184170 75498 184226
rect 75554 184170 75622 184226
rect 75678 184170 85238 184226
rect 85294 184170 85362 184226
rect 85418 184170 93250 184226
rect 93306 184170 93374 184226
rect 93430 184170 93498 184226
rect 93554 184170 93622 184226
rect 93678 184170 111250 184226
rect 111306 184170 111374 184226
rect 111430 184170 111498 184226
rect 111554 184170 111622 184226
rect 111678 184170 115958 184226
rect 116014 184170 116082 184226
rect 116138 184170 146678 184226
rect 146734 184170 146802 184226
rect 146858 184170 177398 184226
rect 177454 184170 177522 184226
rect 177578 184170 208118 184226
rect 208174 184170 208242 184226
rect 208298 184170 238838 184226
rect 238894 184170 238962 184226
rect 239018 184170 269558 184226
rect 269614 184170 269682 184226
rect 269738 184170 300278 184226
rect 300334 184170 300402 184226
rect 300458 184170 330998 184226
rect 331054 184170 331122 184226
rect 331178 184170 361718 184226
rect 361774 184170 361842 184226
rect 361898 184170 392438 184226
rect 392494 184170 392562 184226
rect 392618 184170 423158 184226
rect 423214 184170 423282 184226
rect 423338 184170 453878 184226
rect 453934 184170 454002 184226
rect 454058 184170 484598 184226
rect 484654 184170 484722 184226
rect 484778 184170 515318 184226
rect 515374 184170 515442 184226
rect 515498 184170 546038 184226
rect 546094 184170 546162 184226
rect 546218 184170 561250 184226
rect 561306 184170 561374 184226
rect 561430 184170 561498 184226
rect 561554 184170 561622 184226
rect 561678 184170 579250 184226
rect 579306 184170 579374 184226
rect 579430 184170 579498 184226
rect 579554 184170 579622 184226
rect 579678 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597980 184226
rect -1916 184102 597980 184170
rect -1916 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 3250 184102
rect 3306 184046 3374 184102
rect 3430 184046 3498 184102
rect 3554 184046 3622 184102
rect 3678 184046 21250 184102
rect 21306 184046 21374 184102
rect 21430 184046 21498 184102
rect 21554 184046 21622 184102
rect 21678 184046 39250 184102
rect 39306 184046 39374 184102
rect 39430 184046 39498 184102
rect 39554 184046 39622 184102
rect 39678 184046 54518 184102
rect 54574 184046 54642 184102
rect 54698 184046 57250 184102
rect 57306 184046 57374 184102
rect 57430 184046 57498 184102
rect 57554 184046 57622 184102
rect 57678 184046 75250 184102
rect 75306 184046 75374 184102
rect 75430 184046 75498 184102
rect 75554 184046 75622 184102
rect 75678 184046 85238 184102
rect 85294 184046 85362 184102
rect 85418 184046 93250 184102
rect 93306 184046 93374 184102
rect 93430 184046 93498 184102
rect 93554 184046 93622 184102
rect 93678 184046 111250 184102
rect 111306 184046 111374 184102
rect 111430 184046 111498 184102
rect 111554 184046 111622 184102
rect 111678 184046 115958 184102
rect 116014 184046 116082 184102
rect 116138 184046 146678 184102
rect 146734 184046 146802 184102
rect 146858 184046 177398 184102
rect 177454 184046 177522 184102
rect 177578 184046 208118 184102
rect 208174 184046 208242 184102
rect 208298 184046 238838 184102
rect 238894 184046 238962 184102
rect 239018 184046 269558 184102
rect 269614 184046 269682 184102
rect 269738 184046 300278 184102
rect 300334 184046 300402 184102
rect 300458 184046 330998 184102
rect 331054 184046 331122 184102
rect 331178 184046 361718 184102
rect 361774 184046 361842 184102
rect 361898 184046 392438 184102
rect 392494 184046 392562 184102
rect 392618 184046 423158 184102
rect 423214 184046 423282 184102
rect 423338 184046 453878 184102
rect 453934 184046 454002 184102
rect 454058 184046 484598 184102
rect 484654 184046 484722 184102
rect 484778 184046 515318 184102
rect 515374 184046 515442 184102
rect 515498 184046 546038 184102
rect 546094 184046 546162 184102
rect 546218 184046 561250 184102
rect 561306 184046 561374 184102
rect 561430 184046 561498 184102
rect 561554 184046 561622 184102
rect 561678 184046 579250 184102
rect 579306 184046 579374 184102
rect 579430 184046 579498 184102
rect 579554 184046 579622 184102
rect 579678 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597980 184102
rect -1916 183978 597980 184046
rect -1916 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 3250 183978
rect 3306 183922 3374 183978
rect 3430 183922 3498 183978
rect 3554 183922 3622 183978
rect 3678 183922 21250 183978
rect 21306 183922 21374 183978
rect 21430 183922 21498 183978
rect 21554 183922 21622 183978
rect 21678 183922 39250 183978
rect 39306 183922 39374 183978
rect 39430 183922 39498 183978
rect 39554 183922 39622 183978
rect 39678 183922 54518 183978
rect 54574 183922 54642 183978
rect 54698 183922 57250 183978
rect 57306 183922 57374 183978
rect 57430 183922 57498 183978
rect 57554 183922 57622 183978
rect 57678 183922 75250 183978
rect 75306 183922 75374 183978
rect 75430 183922 75498 183978
rect 75554 183922 75622 183978
rect 75678 183922 85238 183978
rect 85294 183922 85362 183978
rect 85418 183922 93250 183978
rect 93306 183922 93374 183978
rect 93430 183922 93498 183978
rect 93554 183922 93622 183978
rect 93678 183922 111250 183978
rect 111306 183922 111374 183978
rect 111430 183922 111498 183978
rect 111554 183922 111622 183978
rect 111678 183922 115958 183978
rect 116014 183922 116082 183978
rect 116138 183922 146678 183978
rect 146734 183922 146802 183978
rect 146858 183922 177398 183978
rect 177454 183922 177522 183978
rect 177578 183922 208118 183978
rect 208174 183922 208242 183978
rect 208298 183922 238838 183978
rect 238894 183922 238962 183978
rect 239018 183922 269558 183978
rect 269614 183922 269682 183978
rect 269738 183922 300278 183978
rect 300334 183922 300402 183978
rect 300458 183922 330998 183978
rect 331054 183922 331122 183978
rect 331178 183922 361718 183978
rect 361774 183922 361842 183978
rect 361898 183922 392438 183978
rect 392494 183922 392562 183978
rect 392618 183922 423158 183978
rect 423214 183922 423282 183978
rect 423338 183922 453878 183978
rect 453934 183922 454002 183978
rect 454058 183922 484598 183978
rect 484654 183922 484722 183978
rect 484778 183922 515318 183978
rect 515374 183922 515442 183978
rect 515498 183922 546038 183978
rect 546094 183922 546162 183978
rect 546218 183922 561250 183978
rect 561306 183922 561374 183978
rect 561430 183922 561498 183978
rect 561554 183922 561622 183978
rect 561678 183922 579250 183978
rect 579306 183922 579374 183978
rect 579430 183922 579498 183978
rect 579554 183922 579622 183978
rect 579678 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597980 183978
rect -1916 183826 597980 183922
rect -1916 172350 597980 172446
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 6970 172350
rect 7026 172294 7094 172350
rect 7150 172294 7218 172350
rect 7274 172294 7342 172350
rect 7398 172294 24970 172350
rect 25026 172294 25094 172350
rect 25150 172294 25218 172350
rect 25274 172294 25342 172350
rect 25398 172294 42970 172350
rect 43026 172294 43094 172350
rect 43150 172294 43218 172350
rect 43274 172294 43342 172350
rect 43398 172294 60970 172350
rect 61026 172294 61094 172350
rect 61150 172294 61218 172350
rect 61274 172294 61342 172350
rect 61398 172294 69878 172350
rect 69934 172294 70002 172350
rect 70058 172294 78970 172350
rect 79026 172294 79094 172350
rect 79150 172294 79218 172350
rect 79274 172294 79342 172350
rect 79398 172294 96970 172350
rect 97026 172294 97094 172350
rect 97150 172294 97218 172350
rect 97274 172294 97342 172350
rect 97398 172294 100598 172350
rect 100654 172294 100722 172350
rect 100778 172294 131318 172350
rect 131374 172294 131442 172350
rect 131498 172294 162038 172350
rect 162094 172294 162162 172350
rect 162218 172294 192758 172350
rect 192814 172294 192882 172350
rect 192938 172294 223478 172350
rect 223534 172294 223602 172350
rect 223658 172294 254198 172350
rect 254254 172294 254322 172350
rect 254378 172294 284918 172350
rect 284974 172294 285042 172350
rect 285098 172294 315638 172350
rect 315694 172294 315762 172350
rect 315818 172294 346358 172350
rect 346414 172294 346482 172350
rect 346538 172294 377078 172350
rect 377134 172294 377202 172350
rect 377258 172294 407798 172350
rect 407854 172294 407922 172350
rect 407978 172294 438518 172350
rect 438574 172294 438642 172350
rect 438698 172294 469238 172350
rect 469294 172294 469362 172350
rect 469418 172294 499958 172350
rect 500014 172294 500082 172350
rect 500138 172294 530678 172350
rect 530734 172294 530802 172350
rect 530858 172294 564970 172350
rect 565026 172294 565094 172350
rect 565150 172294 565218 172350
rect 565274 172294 565342 172350
rect 565398 172294 582970 172350
rect 583026 172294 583094 172350
rect 583150 172294 583218 172350
rect 583274 172294 583342 172350
rect 583398 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect -1916 172226 597980 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 6970 172226
rect 7026 172170 7094 172226
rect 7150 172170 7218 172226
rect 7274 172170 7342 172226
rect 7398 172170 24970 172226
rect 25026 172170 25094 172226
rect 25150 172170 25218 172226
rect 25274 172170 25342 172226
rect 25398 172170 42970 172226
rect 43026 172170 43094 172226
rect 43150 172170 43218 172226
rect 43274 172170 43342 172226
rect 43398 172170 60970 172226
rect 61026 172170 61094 172226
rect 61150 172170 61218 172226
rect 61274 172170 61342 172226
rect 61398 172170 69878 172226
rect 69934 172170 70002 172226
rect 70058 172170 78970 172226
rect 79026 172170 79094 172226
rect 79150 172170 79218 172226
rect 79274 172170 79342 172226
rect 79398 172170 96970 172226
rect 97026 172170 97094 172226
rect 97150 172170 97218 172226
rect 97274 172170 97342 172226
rect 97398 172170 100598 172226
rect 100654 172170 100722 172226
rect 100778 172170 131318 172226
rect 131374 172170 131442 172226
rect 131498 172170 162038 172226
rect 162094 172170 162162 172226
rect 162218 172170 192758 172226
rect 192814 172170 192882 172226
rect 192938 172170 223478 172226
rect 223534 172170 223602 172226
rect 223658 172170 254198 172226
rect 254254 172170 254322 172226
rect 254378 172170 284918 172226
rect 284974 172170 285042 172226
rect 285098 172170 315638 172226
rect 315694 172170 315762 172226
rect 315818 172170 346358 172226
rect 346414 172170 346482 172226
rect 346538 172170 377078 172226
rect 377134 172170 377202 172226
rect 377258 172170 407798 172226
rect 407854 172170 407922 172226
rect 407978 172170 438518 172226
rect 438574 172170 438642 172226
rect 438698 172170 469238 172226
rect 469294 172170 469362 172226
rect 469418 172170 499958 172226
rect 500014 172170 500082 172226
rect 500138 172170 530678 172226
rect 530734 172170 530802 172226
rect 530858 172170 564970 172226
rect 565026 172170 565094 172226
rect 565150 172170 565218 172226
rect 565274 172170 565342 172226
rect 565398 172170 582970 172226
rect 583026 172170 583094 172226
rect 583150 172170 583218 172226
rect 583274 172170 583342 172226
rect 583398 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect -1916 172102 597980 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 6970 172102
rect 7026 172046 7094 172102
rect 7150 172046 7218 172102
rect 7274 172046 7342 172102
rect 7398 172046 24970 172102
rect 25026 172046 25094 172102
rect 25150 172046 25218 172102
rect 25274 172046 25342 172102
rect 25398 172046 42970 172102
rect 43026 172046 43094 172102
rect 43150 172046 43218 172102
rect 43274 172046 43342 172102
rect 43398 172046 60970 172102
rect 61026 172046 61094 172102
rect 61150 172046 61218 172102
rect 61274 172046 61342 172102
rect 61398 172046 69878 172102
rect 69934 172046 70002 172102
rect 70058 172046 78970 172102
rect 79026 172046 79094 172102
rect 79150 172046 79218 172102
rect 79274 172046 79342 172102
rect 79398 172046 96970 172102
rect 97026 172046 97094 172102
rect 97150 172046 97218 172102
rect 97274 172046 97342 172102
rect 97398 172046 100598 172102
rect 100654 172046 100722 172102
rect 100778 172046 131318 172102
rect 131374 172046 131442 172102
rect 131498 172046 162038 172102
rect 162094 172046 162162 172102
rect 162218 172046 192758 172102
rect 192814 172046 192882 172102
rect 192938 172046 223478 172102
rect 223534 172046 223602 172102
rect 223658 172046 254198 172102
rect 254254 172046 254322 172102
rect 254378 172046 284918 172102
rect 284974 172046 285042 172102
rect 285098 172046 315638 172102
rect 315694 172046 315762 172102
rect 315818 172046 346358 172102
rect 346414 172046 346482 172102
rect 346538 172046 377078 172102
rect 377134 172046 377202 172102
rect 377258 172046 407798 172102
rect 407854 172046 407922 172102
rect 407978 172046 438518 172102
rect 438574 172046 438642 172102
rect 438698 172046 469238 172102
rect 469294 172046 469362 172102
rect 469418 172046 499958 172102
rect 500014 172046 500082 172102
rect 500138 172046 530678 172102
rect 530734 172046 530802 172102
rect 530858 172046 564970 172102
rect 565026 172046 565094 172102
rect 565150 172046 565218 172102
rect 565274 172046 565342 172102
rect 565398 172046 582970 172102
rect 583026 172046 583094 172102
rect 583150 172046 583218 172102
rect 583274 172046 583342 172102
rect 583398 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect -1916 171978 597980 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 6970 171978
rect 7026 171922 7094 171978
rect 7150 171922 7218 171978
rect 7274 171922 7342 171978
rect 7398 171922 24970 171978
rect 25026 171922 25094 171978
rect 25150 171922 25218 171978
rect 25274 171922 25342 171978
rect 25398 171922 42970 171978
rect 43026 171922 43094 171978
rect 43150 171922 43218 171978
rect 43274 171922 43342 171978
rect 43398 171922 60970 171978
rect 61026 171922 61094 171978
rect 61150 171922 61218 171978
rect 61274 171922 61342 171978
rect 61398 171922 69878 171978
rect 69934 171922 70002 171978
rect 70058 171922 78970 171978
rect 79026 171922 79094 171978
rect 79150 171922 79218 171978
rect 79274 171922 79342 171978
rect 79398 171922 96970 171978
rect 97026 171922 97094 171978
rect 97150 171922 97218 171978
rect 97274 171922 97342 171978
rect 97398 171922 100598 171978
rect 100654 171922 100722 171978
rect 100778 171922 131318 171978
rect 131374 171922 131442 171978
rect 131498 171922 162038 171978
rect 162094 171922 162162 171978
rect 162218 171922 192758 171978
rect 192814 171922 192882 171978
rect 192938 171922 223478 171978
rect 223534 171922 223602 171978
rect 223658 171922 254198 171978
rect 254254 171922 254322 171978
rect 254378 171922 284918 171978
rect 284974 171922 285042 171978
rect 285098 171922 315638 171978
rect 315694 171922 315762 171978
rect 315818 171922 346358 171978
rect 346414 171922 346482 171978
rect 346538 171922 377078 171978
rect 377134 171922 377202 171978
rect 377258 171922 407798 171978
rect 407854 171922 407922 171978
rect 407978 171922 438518 171978
rect 438574 171922 438642 171978
rect 438698 171922 469238 171978
rect 469294 171922 469362 171978
rect 469418 171922 499958 171978
rect 500014 171922 500082 171978
rect 500138 171922 530678 171978
rect 530734 171922 530802 171978
rect 530858 171922 564970 171978
rect 565026 171922 565094 171978
rect 565150 171922 565218 171978
rect 565274 171922 565342 171978
rect 565398 171922 582970 171978
rect 583026 171922 583094 171978
rect 583150 171922 583218 171978
rect 583274 171922 583342 171978
rect 583398 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect -1916 171826 597980 171922
rect -1916 166350 597980 166446
rect -1916 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 3250 166350
rect 3306 166294 3374 166350
rect 3430 166294 3498 166350
rect 3554 166294 3622 166350
rect 3678 166294 21250 166350
rect 21306 166294 21374 166350
rect 21430 166294 21498 166350
rect 21554 166294 21622 166350
rect 21678 166294 39250 166350
rect 39306 166294 39374 166350
rect 39430 166294 39498 166350
rect 39554 166294 39622 166350
rect 39678 166294 54518 166350
rect 54574 166294 54642 166350
rect 54698 166294 57250 166350
rect 57306 166294 57374 166350
rect 57430 166294 57498 166350
rect 57554 166294 57622 166350
rect 57678 166294 75250 166350
rect 75306 166294 75374 166350
rect 75430 166294 75498 166350
rect 75554 166294 75622 166350
rect 75678 166294 85238 166350
rect 85294 166294 85362 166350
rect 85418 166294 93250 166350
rect 93306 166294 93374 166350
rect 93430 166294 93498 166350
rect 93554 166294 93622 166350
rect 93678 166294 111250 166350
rect 111306 166294 111374 166350
rect 111430 166294 111498 166350
rect 111554 166294 111622 166350
rect 111678 166294 115958 166350
rect 116014 166294 116082 166350
rect 116138 166294 146678 166350
rect 146734 166294 146802 166350
rect 146858 166294 177398 166350
rect 177454 166294 177522 166350
rect 177578 166294 208118 166350
rect 208174 166294 208242 166350
rect 208298 166294 238838 166350
rect 238894 166294 238962 166350
rect 239018 166294 269558 166350
rect 269614 166294 269682 166350
rect 269738 166294 300278 166350
rect 300334 166294 300402 166350
rect 300458 166294 330998 166350
rect 331054 166294 331122 166350
rect 331178 166294 361718 166350
rect 361774 166294 361842 166350
rect 361898 166294 392438 166350
rect 392494 166294 392562 166350
rect 392618 166294 423158 166350
rect 423214 166294 423282 166350
rect 423338 166294 453878 166350
rect 453934 166294 454002 166350
rect 454058 166294 484598 166350
rect 484654 166294 484722 166350
rect 484778 166294 515318 166350
rect 515374 166294 515442 166350
rect 515498 166294 546038 166350
rect 546094 166294 546162 166350
rect 546218 166294 561250 166350
rect 561306 166294 561374 166350
rect 561430 166294 561498 166350
rect 561554 166294 561622 166350
rect 561678 166294 579250 166350
rect 579306 166294 579374 166350
rect 579430 166294 579498 166350
rect 579554 166294 579622 166350
rect 579678 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597980 166350
rect -1916 166226 597980 166294
rect -1916 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 3250 166226
rect 3306 166170 3374 166226
rect 3430 166170 3498 166226
rect 3554 166170 3622 166226
rect 3678 166170 21250 166226
rect 21306 166170 21374 166226
rect 21430 166170 21498 166226
rect 21554 166170 21622 166226
rect 21678 166170 39250 166226
rect 39306 166170 39374 166226
rect 39430 166170 39498 166226
rect 39554 166170 39622 166226
rect 39678 166170 54518 166226
rect 54574 166170 54642 166226
rect 54698 166170 57250 166226
rect 57306 166170 57374 166226
rect 57430 166170 57498 166226
rect 57554 166170 57622 166226
rect 57678 166170 75250 166226
rect 75306 166170 75374 166226
rect 75430 166170 75498 166226
rect 75554 166170 75622 166226
rect 75678 166170 85238 166226
rect 85294 166170 85362 166226
rect 85418 166170 93250 166226
rect 93306 166170 93374 166226
rect 93430 166170 93498 166226
rect 93554 166170 93622 166226
rect 93678 166170 111250 166226
rect 111306 166170 111374 166226
rect 111430 166170 111498 166226
rect 111554 166170 111622 166226
rect 111678 166170 115958 166226
rect 116014 166170 116082 166226
rect 116138 166170 146678 166226
rect 146734 166170 146802 166226
rect 146858 166170 177398 166226
rect 177454 166170 177522 166226
rect 177578 166170 208118 166226
rect 208174 166170 208242 166226
rect 208298 166170 238838 166226
rect 238894 166170 238962 166226
rect 239018 166170 269558 166226
rect 269614 166170 269682 166226
rect 269738 166170 300278 166226
rect 300334 166170 300402 166226
rect 300458 166170 330998 166226
rect 331054 166170 331122 166226
rect 331178 166170 361718 166226
rect 361774 166170 361842 166226
rect 361898 166170 392438 166226
rect 392494 166170 392562 166226
rect 392618 166170 423158 166226
rect 423214 166170 423282 166226
rect 423338 166170 453878 166226
rect 453934 166170 454002 166226
rect 454058 166170 484598 166226
rect 484654 166170 484722 166226
rect 484778 166170 515318 166226
rect 515374 166170 515442 166226
rect 515498 166170 546038 166226
rect 546094 166170 546162 166226
rect 546218 166170 561250 166226
rect 561306 166170 561374 166226
rect 561430 166170 561498 166226
rect 561554 166170 561622 166226
rect 561678 166170 579250 166226
rect 579306 166170 579374 166226
rect 579430 166170 579498 166226
rect 579554 166170 579622 166226
rect 579678 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597980 166226
rect -1916 166102 597980 166170
rect -1916 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 3250 166102
rect 3306 166046 3374 166102
rect 3430 166046 3498 166102
rect 3554 166046 3622 166102
rect 3678 166046 21250 166102
rect 21306 166046 21374 166102
rect 21430 166046 21498 166102
rect 21554 166046 21622 166102
rect 21678 166046 39250 166102
rect 39306 166046 39374 166102
rect 39430 166046 39498 166102
rect 39554 166046 39622 166102
rect 39678 166046 54518 166102
rect 54574 166046 54642 166102
rect 54698 166046 57250 166102
rect 57306 166046 57374 166102
rect 57430 166046 57498 166102
rect 57554 166046 57622 166102
rect 57678 166046 75250 166102
rect 75306 166046 75374 166102
rect 75430 166046 75498 166102
rect 75554 166046 75622 166102
rect 75678 166046 85238 166102
rect 85294 166046 85362 166102
rect 85418 166046 93250 166102
rect 93306 166046 93374 166102
rect 93430 166046 93498 166102
rect 93554 166046 93622 166102
rect 93678 166046 111250 166102
rect 111306 166046 111374 166102
rect 111430 166046 111498 166102
rect 111554 166046 111622 166102
rect 111678 166046 115958 166102
rect 116014 166046 116082 166102
rect 116138 166046 146678 166102
rect 146734 166046 146802 166102
rect 146858 166046 177398 166102
rect 177454 166046 177522 166102
rect 177578 166046 208118 166102
rect 208174 166046 208242 166102
rect 208298 166046 238838 166102
rect 238894 166046 238962 166102
rect 239018 166046 269558 166102
rect 269614 166046 269682 166102
rect 269738 166046 300278 166102
rect 300334 166046 300402 166102
rect 300458 166046 330998 166102
rect 331054 166046 331122 166102
rect 331178 166046 361718 166102
rect 361774 166046 361842 166102
rect 361898 166046 392438 166102
rect 392494 166046 392562 166102
rect 392618 166046 423158 166102
rect 423214 166046 423282 166102
rect 423338 166046 453878 166102
rect 453934 166046 454002 166102
rect 454058 166046 484598 166102
rect 484654 166046 484722 166102
rect 484778 166046 515318 166102
rect 515374 166046 515442 166102
rect 515498 166046 546038 166102
rect 546094 166046 546162 166102
rect 546218 166046 561250 166102
rect 561306 166046 561374 166102
rect 561430 166046 561498 166102
rect 561554 166046 561622 166102
rect 561678 166046 579250 166102
rect 579306 166046 579374 166102
rect 579430 166046 579498 166102
rect 579554 166046 579622 166102
rect 579678 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597980 166102
rect -1916 165978 597980 166046
rect -1916 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 3250 165978
rect 3306 165922 3374 165978
rect 3430 165922 3498 165978
rect 3554 165922 3622 165978
rect 3678 165922 21250 165978
rect 21306 165922 21374 165978
rect 21430 165922 21498 165978
rect 21554 165922 21622 165978
rect 21678 165922 39250 165978
rect 39306 165922 39374 165978
rect 39430 165922 39498 165978
rect 39554 165922 39622 165978
rect 39678 165922 54518 165978
rect 54574 165922 54642 165978
rect 54698 165922 57250 165978
rect 57306 165922 57374 165978
rect 57430 165922 57498 165978
rect 57554 165922 57622 165978
rect 57678 165922 75250 165978
rect 75306 165922 75374 165978
rect 75430 165922 75498 165978
rect 75554 165922 75622 165978
rect 75678 165922 85238 165978
rect 85294 165922 85362 165978
rect 85418 165922 93250 165978
rect 93306 165922 93374 165978
rect 93430 165922 93498 165978
rect 93554 165922 93622 165978
rect 93678 165922 111250 165978
rect 111306 165922 111374 165978
rect 111430 165922 111498 165978
rect 111554 165922 111622 165978
rect 111678 165922 115958 165978
rect 116014 165922 116082 165978
rect 116138 165922 146678 165978
rect 146734 165922 146802 165978
rect 146858 165922 177398 165978
rect 177454 165922 177522 165978
rect 177578 165922 208118 165978
rect 208174 165922 208242 165978
rect 208298 165922 238838 165978
rect 238894 165922 238962 165978
rect 239018 165922 269558 165978
rect 269614 165922 269682 165978
rect 269738 165922 300278 165978
rect 300334 165922 300402 165978
rect 300458 165922 330998 165978
rect 331054 165922 331122 165978
rect 331178 165922 361718 165978
rect 361774 165922 361842 165978
rect 361898 165922 392438 165978
rect 392494 165922 392562 165978
rect 392618 165922 423158 165978
rect 423214 165922 423282 165978
rect 423338 165922 453878 165978
rect 453934 165922 454002 165978
rect 454058 165922 484598 165978
rect 484654 165922 484722 165978
rect 484778 165922 515318 165978
rect 515374 165922 515442 165978
rect 515498 165922 546038 165978
rect 546094 165922 546162 165978
rect 546218 165922 561250 165978
rect 561306 165922 561374 165978
rect 561430 165922 561498 165978
rect 561554 165922 561622 165978
rect 561678 165922 579250 165978
rect 579306 165922 579374 165978
rect 579430 165922 579498 165978
rect 579554 165922 579622 165978
rect 579678 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597980 165978
rect -1916 165826 597980 165922
rect -1916 154350 597980 154446
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 6970 154350
rect 7026 154294 7094 154350
rect 7150 154294 7218 154350
rect 7274 154294 7342 154350
rect 7398 154294 24970 154350
rect 25026 154294 25094 154350
rect 25150 154294 25218 154350
rect 25274 154294 25342 154350
rect 25398 154294 42970 154350
rect 43026 154294 43094 154350
rect 43150 154294 43218 154350
rect 43274 154294 43342 154350
rect 43398 154294 60970 154350
rect 61026 154294 61094 154350
rect 61150 154294 61218 154350
rect 61274 154294 61342 154350
rect 61398 154294 69878 154350
rect 69934 154294 70002 154350
rect 70058 154294 78970 154350
rect 79026 154294 79094 154350
rect 79150 154294 79218 154350
rect 79274 154294 79342 154350
rect 79398 154294 96970 154350
rect 97026 154294 97094 154350
rect 97150 154294 97218 154350
rect 97274 154294 97342 154350
rect 97398 154294 100598 154350
rect 100654 154294 100722 154350
rect 100778 154294 131318 154350
rect 131374 154294 131442 154350
rect 131498 154294 162038 154350
rect 162094 154294 162162 154350
rect 162218 154294 192758 154350
rect 192814 154294 192882 154350
rect 192938 154294 223478 154350
rect 223534 154294 223602 154350
rect 223658 154294 254198 154350
rect 254254 154294 254322 154350
rect 254378 154294 284918 154350
rect 284974 154294 285042 154350
rect 285098 154294 315638 154350
rect 315694 154294 315762 154350
rect 315818 154294 346358 154350
rect 346414 154294 346482 154350
rect 346538 154294 377078 154350
rect 377134 154294 377202 154350
rect 377258 154294 407798 154350
rect 407854 154294 407922 154350
rect 407978 154294 438518 154350
rect 438574 154294 438642 154350
rect 438698 154294 469238 154350
rect 469294 154294 469362 154350
rect 469418 154294 499958 154350
rect 500014 154294 500082 154350
rect 500138 154294 530678 154350
rect 530734 154294 530802 154350
rect 530858 154294 564970 154350
rect 565026 154294 565094 154350
rect 565150 154294 565218 154350
rect 565274 154294 565342 154350
rect 565398 154294 582970 154350
rect 583026 154294 583094 154350
rect 583150 154294 583218 154350
rect 583274 154294 583342 154350
rect 583398 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect -1916 154226 597980 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 6970 154226
rect 7026 154170 7094 154226
rect 7150 154170 7218 154226
rect 7274 154170 7342 154226
rect 7398 154170 24970 154226
rect 25026 154170 25094 154226
rect 25150 154170 25218 154226
rect 25274 154170 25342 154226
rect 25398 154170 42970 154226
rect 43026 154170 43094 154226
rect 43150 154170 43218 154226
rect 43274 154170 43342 154226
rect 43398 154170 60970 154226
rect 61026 154170 61094 154226
rect 61150 154170 61218 154226
rect 61274 154170 61342 154226
rect 61398 154170 69878 154226
rect 69934 154170 70002 154226
rect 70058 154170 78970 154226
rect 79026 154170 79094 154226
rect 79150 154170 79218 154226
rect 79274 154170 79342 154226
rect 79398 154170 96970 154226
rect 97026 154170 97094 154226
rect 97150 154170 97218 154226
rect 97274 154170 97342 154226
rect 97398 154170 100598 154226
rect 100654 154170 100722 154226
rect 100778 154170 131318 154226
rect 131374 154170 131442 154226
rect 131498 154170 162038 154226
rect 162094 154170 162162 154226
rect 162218 154170 192758 154226
rect 192814 154170 192882 154226
rect 192938 154170 223478 154226
rect 223534 154170 223602 154226
rect 223658 154170 254198 154226
rect 254254 154170 254322 154226
rect 254378 154170 284918 154226
rect 284974 154170 285042 154226
rect 285098 154170 315638 154226
rect 315694 154170 315762 154226
rect 315818 154170 346358 154226
rect 346414 154170 346482 154226
rect 346538 154170 377078 154226
rect 377134 154170 377202 154226
rect 377258 154170 407798 154226
rect 407854 154170 407922 154226
rect 407978 154170 438518 154226
rect 438574 154170 438642 154226
rect 438698 154170 469238 154226
rect 469294 154170 469362 154226
rect 469418 154170 499958 154226
rect 500014 154170 500082 154226
rect 500138 154170 530678 154226
rect 530734 154170 530802 154226
rect 530858 154170 564970 154226
rect 565026 154170 565094 154226
rect 565150 154170 565218 154226
rect 565274 154170 565342 154226
rect 565398 154170 582970 154226
rect 583026 154170 583094 154226
rect 583150 154170 583218 154226
rect 583274 154170 583342 154226
rect 583398 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect -1916 154102 597980 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 6970 154102
rect 7026 154046 7094 154102
rect 7150 154046 7218 154102
rect 7274 154046 7342 154102
rect 7398 154046 24970 154102
rect 25026 154046 25094 154102
rect 25150 154046 25218 154102
rect 25274 154046 25342 154102
rect 25398 154046 42970 154102
rect 43026 154046 43094 154102
rect 43150 154046 43218 154102
rect 43274 154046 43342 154102
rect 43398 154046 60970 154102
rect 61026 154046 61094 154102
rect 61150 154046 61218 154102
rect 61274 154046 61342 154102
rect 61398 154046 69878 154102
rect 69934 154046 70002 154102
rect 70058 154046 78970 154102
rect 79026 154046 79094 154102
rect 79150 154046 79218 154102
rect 79274 154046 79342 154102
rect 79398 154046 96970 154102
rect 97026 154046 97094 154102
rect 97150 154046 97218 154102
rect 97274 154046 97342 154102
rect 97398 154046 100598 154102
rect 100654 154046 100722 154102
rect 100778 154046 131318 154102
rect 131374 154046 131442 154102
rect 131498 154046 162038 154102
rect 162094 154046 162162 154102
rect 162218 154046 192758 154102
rect 192814 154046 192882 154102
rect 192938 154046 223478 154102
rect 223534 154046 223602 154102
rect 223658 154046 254198 154102
rect 254254 154046 254322 154102
rect 254378 154046 284918 154102
rect 284974 154046 285042 154102
rect 285098 154046 315638 154102
rect 315694 154046 315762 154102
rect 315818 154046 346358 154102
rect 346414 154046 346482 154102
rect 346538 154046 377078 154102
rect 377134 154046 377202 154102
rect 377258 154046 407798 154102
rect 407854 154046 407922 154102
rect 407978 154046 438518 154102
rect 438574 154046 438642 154102
rect 438698 154046 469238 154102
rect 469294 154046 469362 154102
rect 469418 154046 499958 154102
rect 500014 154046 500082 154102
rect 500138 154046 530678 154102
rect 530734 154046 530802 154102
rect 530858 154046 564970 154102
rect 565026 154046 565094 154102
rect 565150 154046 565218 154102
rect 565274 154046 565342 154102
rect 565398 154046 582970 154102
rect 583026 154046 583094 154102
rect 583150 154046 583218 154102
rect 583274 154046 583342 154102
rect 583398 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect -1916 153978 597980 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 6970 153978
rect 7026 153922 7094 153978
rect 7150 153922 7218 153978
rect 7274 153922 7342 153978
rect 7398 153922 24970 153978
rect 25026 153922 25094 153978
rect 25150 153922 25218 153978
rect 25274 153922 25342 153978
rect 25398 153922 42970 153978
rect 43026 153922 43094 153978
rect 43150 153922 43218 153978
rect 43274 153922 43342 153978
rect 43398 153922 60970 153978
rect 61026 153922 61094 153978
rect 61150 153922 61218 153978
rect 61274 153922 61342 153978
rect 61398 153922 69878 153978
rect 69934 153922 70002 153978
rect 70058 153922 78970 153978
rect 79026 153922 79094 153978
rect 79150 153922 79218 153978
rect 79274 153922 79342 153978
rect 79398 153922 96970 153978
rect 97026 153922 97094 153978
rect 97150 153922 97218 153978
rect 97274 153922 97342 153978
rect 97398 153922 100598 153978
rect 100654 153922 100722 153978
rect 100778 153922 131318 153978
rect 131374 153922 131442 153978
rect 131498 153922 162038 153978
rect 162094 153922 162162 153978
rect 162218 153922 192758 153978
rect 192814 153922 192882 153978
rect 192938 153922 223478 153978
rect 223534 153922 223602 153978
rect 223658 153922 254198 153978
rect 254254 153922 254322 153978
rect 254378 153922 284918 153978
rect 284974 153922 285042 153978
rect 285098 153922 315638 153978
rect 315694 153922 315762 153978
rect 315818 153922 346358 153978
rect 346414 153922 346482 153978
rect 346538 153922 377078 153978
rect 377134 153922 377202 153978
rect 377258 153922 407798 153978
rect 407854 153922 407922 153978
rect 407978 153922 438518 153978
rect 438574 153922 438642 153978
rect 438698 153922 469238 153978
rect 469294 153922 469362 153978
rect 469418 153922 499958 153978
rect 500014 153922 500082 153978
rect 500138 153922 530678 153978
rect 530734 153922 530802 153978
rect 530858 153922 564970 153978
rect 565026 153922 565094 153978
rect 565150 153922 565218 153978
rect 565274 153922 565342 153978
rect 565398 153922 582970 153978
rect 583026 153922 583094 153978
rect 583150 153922 583218 153978
rect 583274 153922 583342 153978
rect 583398 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect -1916 153826 597980 153922
rect -1916 148350 597980 148446
rect -1916 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 3250 148350
rect 3306 148294 3374 148350
rect 3430 148294 3498 148350
rect 3554 148294 3622 148350
rect 3678 148294 21250 148350
rect 21306 148294 21374 148350
rect 21430 148294 21498 148350
rect 21554 148294 21622 148350
rect 21678 148294 39250 148350
rect 39306 148294 39374 148350
rect 39430 148294 39498 148350
rect 39554 148294 39622 148350
rect 39678 148294 54518 148350
rect 54574 148294 54642 148350
rect 54698 148294 57250 148350
rect 57306 148294 57374 148350
rect 57430 148294 57498 148350
rect 57554 148294 57622 148350
rect 57678 148294 75250 148350
rect 75306 148294 75374 148350
rect 75430 148294 75498 148350
rect 75554 148294 75622 148350
rect 75678 148294 85238 148350
rect 85294 148294 85362 148350
rect 85418 148294 93250 148350
rect 93306 148294 93374 148350
rect 93430 148294 93498 148350
rect 93554 148294 93622 148350
rect 93678 148294 111250 148350
rect 111306 148294 111374 148350
rect 111430 148294 111498 148350
rect 111554 148294 111622 148350
rect 111678 148294 115958 148350
rect 116014 148294 116082 148350
rect 116138 148294 146678 148350
rect 146734 148294 146802 148350
rect 146858 148294 177398 148350
rect 177454 148294 177522 148350
rect 177578 148294 208118 148350
rect 208174 148294 208242 148350
rect 208298 148294 238838 148350
rect 238894 148294 238962 148350
rect 239018 148294 269558 148350
rect 269614 148294 269682 148350
rect 269738 148294 300278 148350
rect 300334 148294 300402 148350
rect 300458 148294 330998 148350
rect 331054 148294 331122 148350
rect 331178 148294 361718 148350
rect 361774 148294 361842 148350
rect 361898 148294 392438 148350
rect 392494 148294 392562 148350
rect 392618 148294 423158 148350
rect 423214 148294 423282 148350
rect 423338 148294 453878 148350
rect 453934 148294 454002 148350
rect 454058 148294 484598 148350
rect 484654 148294 484722 148350
rect 484778 148294 515318 148350
rect 515374 148294 515442 148350
rect 515498 148294 546038 148350
rect 546094 148294 546162 148350
rect 546218 148294 561250 148350
rect 561306 148294 561374 148350
rect 561430 148294 561498 148350
rect 561554 148294 561622 148350
rect 561678 148294 579250 148350
rect 579306 148294 579374 148350
rect 579430 148294 579498 148350
rect 579554 148294 579622 148350
rect 579678 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597980 148350
rect -1916 148226 597980 148294
rect -1916 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 3250 148226
rect 3306 148170 3374 148226
rect 3430 148170 3498 148226
rect 3554 148170 3622 148226
rect 3678 148170 21250 148226
rect 21306 148170 21374 148226
rect 21430 148170 21498 148226
rect 21554 148170 21622 148226
rect 21678 148170 39250 148226
rect 39306 148170 39374 148226
rect 39430 148170 39498 148226
rect 39554 148170 39622 148226
rect 39678 148170 54518 148226
rect 54574 148170 54642 148226
rect 54698 148170 57250 148226
rect 57306 148170 57374 148226
rect 57430 148170 57498 148226
rect 57554 148170 57622 148226
rect 57678 148170 75250 148226
rect 75306 148170 75374 148226
rect 75430 148170 75498 148226
rect 75554 148170 75622 148226
rect 75678 148170 85238 148226
rect 85294 148170 85362 148226
rect 85418 148170 93250 148226
rect 93306 148170 93374 148226
rect 93430 148170 93498 148226
rect 93554 148170 93622 148226
rect 93678 148170 111250 148226
rect 111306 148170 111374 148226
rect 111430 148170 111498 148226
rect 111554 148170 111622 148226
rect 111678 148170 115958 148226
rect 116014 148170 116082 148226
rect 116138 148170 146678 148226
rect 146734 148170 146802 148226
rect 146858 148170 177398 148226
rect 177454 148170 177522 148226
rect 177578 148170 208118 148226
rect 208174 148170 208242 148226
rect 208298 148170 238838 148226
rect 238894 148170 238962 148226
rect 239018 148170 269558 148226
rect 269614 148170 269682 148226
rect 269738 148170 300278 148226
rect 300334 148170 300402 148226
rect 300458 148170 330998 148226
rect 331054 148170 331122 148226
rect 331178 148170 361718 148226
rect 361774 148170 361842 148226
rect 361898 148170 392438 148226
rect 392494 148170 392562 148226
rect 392618 148170 423158 148226
rect 423214 148170 423282 148226
rect 423338 148170 453878 148226
rect 453934 148170 454002 148226
rect 454058 148170 484598 148226
rect 484654 148170 484722 148226
rect 484778 148170 515318 148226
rect 515374 148170 515442 148226
rect 515498 148170 546038 148226
rect 546094 148170 546162 148226
rect 546218 148170 561250 148226
rect 561306 148170 561374 148226
rect 561430 148170 561498 148226
rect 561554 148170 561622 148226
rect 561678 148170 579250 148226
rect 579306 148170 579374 148226
rect 579430 148170 579498 148226
rect 579554 148170 579622 148226
rect 579678 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597980 148226
rect -1916 148102 597980 148170
rect -1916 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 3250 148102
rect 3306 148046 3374 148102
rect 3430 148046 3498 148102
rect 3554 148046 3622 148102
rect 3678 148046 21250 148102
rect 21306 148046 21374 148102
rect 21430 148046 21498 148102
rect 21554 148046 21622 148102
rect 21678 148046 39250 148102
rect 39306 148046 39374 148102
rect 39430 148046 39498 148102
rect 39554 148046 39622 148102
rect 39678 148046 54518 148102
rect 54574 148046 54642 148102
rect 54698 148046 57250 148102
rect 57306 148046 57374 148102
rect 57430 148046 57498 148102
rect 57554 148046 57622 148102
rect 57678 148046 75250 148102
rect 75306 148046 75374 148102
rect 75430 148046 75498 148102
rect 75554 148046 75622 148102
rect 75678 148046 85238 148102
rect 85294 148046 85362 148102
rect 85418 148046 93250 148102
rect 93306 148046 93374 148102
rect 93430 148046 93498 148102
rect 93554 148046 93622 148102
rect 93678 148046 111250 148102
rect 111306 148046 111374 148102
rect 111430 148046 111498 148102
rect 111554 148046 111622 148102
rect 111678 148046 115958 148102
rect 116014 148046 116082 148102
rect 116138 148046 146678 148102
rect 146734 148046 146802 148102
rect 146858 148046 177398 148102
rect 177454 148046 177522 148102
rect 177578 148046 208118 148102
rect 208174 148046 208242 148102
rect 208298 148046 238838 148102
rect 238894 148046 238962 148102
rect 239018 148046 269558 148102
rect 269614 148046 269682 148102
rect 269738 148046 300278 148102
rect 300334 148046 300402 148102
rect 300458 148046 330998 148102
rect 331054 148046 331122 148102
rect 331178 148046 361718 148102
rect 361774 148046 361842 148102
rect 361898 148046 392438 148102
rect 392494 148046 392562 148102
rect 392618 148046 423158 148102
rect 423214 148046 423282 148102
rect 423338 148046 453878 148102
rect 453934 148046 454002 148102
rect 454058 148046 484598 148102
rect 484654 148046 484722 148102
rect 484778 148046 515318 148102
rect 515374 148046 515442 148102
rect 515498 148046 546038 148102
rect 546094 148046 546162 148102
rect 546218 148046 561250 148102
rect 561306 148046 561374 148102
rect 561430 148046 561498 148102
rect 561554 148046 561622 148102
rect 561678 148046 579250 148102
rect 579306 148046 579374 148102
rect 579430 148046 579498 148102
rect 579554 148046 579622 148102
rect 579678 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597980 148102
rect -1916 147978 597980 148046
rect -1916 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 3250 147978
rect 3306 147922 3374 147978
rect 3430 147922 3498 147978
rect 3554 147922 3622 147978
rect 3678 147922 21250 147978
rect 21306 147922 21374 147978
rect 21430 147922 21498 147978
rect 21554 147922 21622 147978
rect 21678 147922 39250 147978
rect 39306 147922 39374 147978
rect 39430 147922 39498 147978
rect 39554 147922 39622 147978
rect 39678 147922 54518 147978
rect 54574 147922 54642 147978
rect 54698 147922 57250 147978
rect 57306 147922 57374 147978
rect 57430 147922 57498 147978
rect 57554 147922 57622 147978
rect 57678 147922 75250 147978
rect 75306 147922 75374 147978
rect 75430 147922 75498 147978
rect 75554 147922 75622 147978
rect 75678 147922 85238 147978
rect 85294 147922 85362 147978
rect 85418 147922 93250 147978
rect 93306 147922 93374 147978
rect 93430 147922 93498 147978
rect 93554 147922 93622 147978
rect 93678 147922 111250 147978
rect 111306 147922 111374 147978
rect 111430 147922 111498 147978
rect 111554 147922 111622 147978
rect 111678 147922 115958 147978
rect 116014 147922 116082 147978
rect 116138 147922 146678 147978
rect 146734 147922 146802 147978
rect 146858 147922 177398 147978
rect 177454 147922 177522 147978
rect 177578 147922 208118 147978
rect 208174 147922 208242 147978
rect 208298 147922 238838 147978
rect 238894 147922 238962 147978
rect 239018 147922 269558 147978
rect 269614 147922 269682 147978
rect 269738 147922 300278 147978
rect 300334 147922 300402 147978
rect 300458 147922 330998 147978
rect 331054 147922 331122 147978
rect 331178 147922 361718 147978
rect 361774 147922 361842 147978
rect 361898 147922 392438 147978
rect 392494 147922 392562 147978
rect 392618 147922 423158 147978
rect 423214 147922 423282 147978
rect 423338 147922 453878 147978
rect 453934 147922 454002 147978
rect 454058 147922 484598 147978
rect 484654 147922 484722 147978
rect 484778 147922 515318 147978
rect 515374 147922 515442 147978
rect 515498 147922 546038 147978
rect 546094 147922 546162 147978
rect 546218 147922 561250 147978
rect 561306 147922 561374 147978
rect 561430 147922 561498 147978
rect 561554 147922 561622 147978
rect 561678 147922 579250 147978
rect 579306 147922 579374 147978
rect 579430 147922 579498 147978
rect 579554 147922 579622 147978
rect 579678 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597980 147978
rect -1916 147826 597980 147922
rect -1916 136350 597980 136446
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 6970 136350
rect 7026 136294 7094 136350
rect 7150 136294 7218 136350
rect 7274 136294 7342 136350
rect 7398 136294 24970 136350
rect 25026 136294 25094 136350
rect 25150 136294 25218 136350
rect 25274 136294 25342 136350
rect 25398 136294 42970 136350
rect 43026 136294 43094 136350
rect 43150 136294 43218 136350
rect 43274 136294 43342 136350
rect 43398 136294 60970 136350
rect 61026 136294 61094 136350
rect 61150 136294 61218 136350
rect 61274 136294 61342 136350
rect 61398 136294 69878 136350
rect 69934 136294 70002 136350
rect 70058 136294 78970 136350
rect 79026 136294 79094 136350
rect 79150 136294 79218 136350
rect 79274 136294 79342 136350
rect 79398 136294 96970 136350
rect 97026 136294 97094 136350
rect 97150 136294 97218 136350
rect 97274 136294 97342 136350
rect 97398 136294 100598 136350
rect 100654 136294 100722 136350
rect 100778 136294 131318 136350
rect 131374 136294 131442 136350
rect 131498 136294 162038 136350
rect 162094 136294 162162 136350
rect 162218 136294 192758 136350
rect 192814 136294 192882 136350
rect 192938 136294 223478 136350
rect 223534 136294 223602 136350
rect 223658 136294 254198 136350
rect 254254 136294 254322 136350
rect 254378 136294 284918 136350
rect 284974 136294 285042 136350
rect 285098 136294 315638 136350
rect 315694 136294 315762 136350
rect 315818 136294 346358 136350
rect 346414 136294 346482 136350
rect 346538 136294 377078 136350
rect 377134 136294 377202 136350
rect 377258 136294 407798 136350
rect 407854 136294 407922 136350
rect 407978 136294 438518 136350
rect 438574 136294 438642 136350
rect 438698 136294 469238 136350
rect 469294 136294 469362 136350
rect 469418 136294 499958 136350
rect 500014 136294 500082 136350
rect 500138 136294 530678 136350
rect 530734 136294 530802 136350
rect 530858 136294 564970 136350
rect 565026 136294 565094 136350
rect 565150 136294 565218 136350
rect 565274 136294 565342 136350
rect 565398 136294 582970 136350
rect 583026 136294 583094 136350
rect 583150 136294 583218 136350
rect 583274 136294 583342 136350
rect 583398 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect -1916 136226 597980 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 6970 136226
rect 7026 136170 7094 136226
rect 7150 136170 7218 136226
rect 7274 136170 7342 136226
rect 7398 136170 24970 136226
rect 25026 136170 25094 136226
rect 25150 136170 25218 136226
rect 25274 136170 25342 136226
rect 25398 136170 42970 136226
rect 43026 136170 43094 136226
rect 43150 136170 43218 136226
rect 43274 136170 43342 136226
rect 43398 136170 60970 136226
rect 61026 136170 61094 136226
rect 61150 136170 61218 136226
rect 61274 136170 61342 136226
rect 61398 136170 69878 136226
rect 69934 136170 70002 136226
rect 70058 136170 78970 136226
rect 79026 136170 79094 136226
rect 79150 136170 79218 136226
rect 79274 136170 79342 136226
rect 79398 136170 96970 136226
rect 97026 136170 97094 136226
rect 97150 136170 97218 136226
rect 97274 136170 97342 136226
rect 97398 136170 100598 136226
rect 100654 136170 100722 136226
rect 100778 136170 131318 136226
rect 131374 136170 131442 136226
rect 131498 136170 162038 136226
rect 162094 136170 162162 136226
rect 162218 136170 192758 136226
rect 192814 136170 192882 136226
rect 192938 136170 223478 136226
rect 223534 136170 223602 136226
rect 223658 136170 254198 136226
rect 254254 136170 254322 136226
rect 254378 136170 284918 136226
rect 284974 136170 285042 136226
rect 285098 136170 315638 136226
rect 315694 136170 315762 136226
rect 315818 136170 346358 136226
rect 346414 136170 346482 136226
rect 346538 136170 377078 136226
rect 377134 136170 377202 136226
rect 377258 136170 407798 136226
rect 407854 136170 407922 136226
rect 407978 136170 438518 136226
rect 438574 136170 438642 136226
rect 438698 136170 469238 136226
rect 469294 136170 469362 136226
rect 469418 136170 499958 136226
rect 500014 136170 500082 136226
rect 500138 136170 530678 136226
rect 530734 136170 530802 136226
rect 530858 136170 564970 136226
rect 565026 136170 565094 136226
rect 565150 136170 565218 136226
rect 565274 136170 565342 136226
rect 565398 136170 582970 136226
rect 583026 136170 583094 136226
rect 583150 136170 583218 136226
rect 583274 136170 583342 136226
rect 583398 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect -1916 136102 597980 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 6970 136102
rect 7026 136046 7094 136102
rect 7150 136046 7218 136102
rect 7274 136046 7342 136102
rect 7398 136046 24970 136102
rect 25026 136046 25094 136102
rect 25150 136046 25218 136102
rect 25274 136046 25342 136102
rect 25398 136046 42970 136102
rect 43026 136046 43094 136102
rect 43150 136046 43218 136102
rect 43274 136046 43342 136102
rect 43398 136046 60970 136102
rect 61026 136046 61094 136102
rect 61150 136046 61218 136102
rect 61274 136046 61342 136102
rect 61398 136046 69878 136102
rect 69934 136046 70002 136102
rect 70058 136046 78970 136102
rect 79026 136046 79094 136102
rect 79150 136046 79218 136102
rect 79274 136046 79342 136102
rect 79398 136046 96970 136102
rect 97026 136046 97094 136102
rect 97150 136046 97218 136102
rect 97274 136046 97342 136102
rect 97398 136046 100598 136102
rect 100654 136046 100722 136102
rect 100778 136046 131318 136102
rect 131374 136046 131442 136102
rect 131498 136046 162038 136102
rect 162094 136046 162162 136102
rect 162218 136046 192758 136102
rect 192814 136046 192882 136102
rect 192938 136046 223478 136102
rect 223534 136046 223602 136102
rect 223658 136046 254198 136102
rect 254254 136046 254322 136102
rect 254378 136046 284918 136102
rect 284974 136046 285042 136102
rect 285098 136046 315638 136102
rect 315694 136046 315762 136102
rect 315818 136046 346358 136102
rect 346414 136046 346482 136102
rect 346538 136046 377078 136102
rect 377134 136046 377202 136102
rect 377258 136046 407798 136102
rect 407854 136046 407922 136102
rect 407978 136046 438518 136102
rect 438574 136046 438642 136102
rect 438698 136046 469238 136102
rect 469294 136046 469362 136102
rect 469418 136046 499958 136102
rect 500014 136046 500082 136102
rect 500138 136046 530678 136102
rect 530734 136046 530802 136102
rect 530858 136046 564970 136102
rect 565026 136046 565094 136102
rect 565150 136046 565218 136102
rect 565274 136046 565342 136102
rect 565398 136046 582970 136102
rect 583026 136046 583094 136102
rect 583150 136046 583218 136102
rect 583274 136046 583342 136102
rect 583398 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect -1916 135978 597980 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 6970 135978
rect 7026 135922 7094 135978
rect 7150 135922 7218 135978
rect 7274 135922 7342 135978
rect 7398 135922 24970 135978
rect 25026 135922 25094 135978
rect 25150 135922 25218 135978
rect 25274 135922 25342 135978
rect 25398 135922 42970 135978
rect 43026 135922 43094 135978
rect 43150 135922 43218 135978
rect 43274 135922 43342 135978
rect 43398 135922 60970 135978
rect 61026 135922 61094 135978
rect 61150 135922 61218 135978
rect 61274 135922 61342 135978
rect 61398 135922 69878 135978
rect 69934 135922 70002 135978
rect 70058 135922 78970 135978
rect 79026 135922 79094 135978
rect 79150 135922 79218 135978
rect 79274 135922 79342 135978
rect 79398 135922 96970 135978
rect 97026 135922 97094 135978
rect 97150 135922 97218 135978
rect 97274 135922 97342 135978
rect 97398 135922 100598 135978
rect 100654 135922 100722 135978
rect 100778 135922 131318 135978
rect 131374 135922 131442 135978
rect 131498 135922 162038 135978
rect 162094 135922 162162 135978
rect 162218 135922 192758 135978
rect 192814 135922 192882 135978
rect 192938 135922 223478 135978
rect 223534 135922 223602 135978
rect 223658 135922 254198 135978
rect 254254 135922 254322 135978
rect 254378 135922 284918 135978
rect 284974 135922 285042 135978
rect 285098 135922 315638 135978
rect 315694 135922 315762 135978
rect 315818 135922 346358 135978
rect 346414 135922 346482 135978
rect 346538 135922 377078 135978
rect 377134 135922 377202 135978
rect 377258 135922 407798 135978
rect 407854 135922 407922 135978
rect 407978 135922 438518 135978
rect 438574 135922 438642 135978
rect 438698 135922 469238 135978
rect 469294 135922 469362 135978
rect 469418 135922 499958 135978
rect 500014 135922 500082 135978
rect 500138 135922 530678 135978
rect 530734 135922 530802 135978
rect 530858 135922 564970 135978
rect 565026 135922 565094 135978
rect 565150 135922 565218 135978
rect 565274 135922 565342 135978
rect 565398 135922 582970 135978
rect 583026 135922 583094 135978
rect 583150 135922 583218 135978
rect 583274 135922 583342 135978
rect 583398 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect -1916 135826 597980 135922
rect -1916 130350 597980 130446
rect -1916 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 3250 130350
rect 3306 130294 3374 130350
rect 3430 130294 3498 130350
rect 3554 130294 3622 130350
rect 3678 130294 21250 130350
rect 21306 130294 21374 130350
rect 21430 130294 21498 130350
rect 21554 130294 21622 130350
rect 21678 130294 39250 130350
rect 39306 130294 39374 130350
rect 39430 130294 39498 130350
rect 39554 130294 39622 130350
rect 39678 130294 54518 130350
rect 54574 130294 54642 130350
rect 54698 130294 57250 130350
rect 57306 130294 57374 130350
rect 57430 130294 57498 130350
rect 57554 130294 57622 130350
rect 57678 130294 75250 130350
rect 75306 130294 75374 130350
rect 75430 130294 75498 130350
rect 75554 130294 75622 130350
rect 75678 130294 85238 130350
rect 85294 130294 85362 130350
rect 85418 130294 93250 130350
rect 93306 130294 93374 130350
rect 93430 130294 93498 130350
rect 93554 130294 93622 130350
rect 93678 130294 111250 130350
rect 111306 130294 111374 130350
rect 111430 130294 111498 130350
rect 111554 130294 111622 130350
rect 111678 130294 115958 130350
rect 116014 130294 116082 130350
rect 116138 130294 146678 130350
rect 146734 130294 146802 130350
rect 146858 130294 177398 130350
rect 177454 130294 177522 130350
rect 177578 130294 208118 130350
rect 208174 130294 208242 130350
rect 208298 130294 238838 130350
rect 238894 130294 238962 130350
rect 239018 130294 269558 130350
rect 269614 130294 269682 130350
rect 269738 130294 300278 130350
rect 300334 130294 300402 130350
rect 300458 130294 330998 130350
rect 331054 130294 331122 130350
rect 331178 130294 361718 130350
rect 361774 130294 361842 130350
rect 361898 130294 392438 130350
rect 392494 130294 392562 130350
rect 392618 130294 423158 130350
rect 423214 130294 423282 130350
rect 423338 130294 453878 130350
rect 453934 130294 454002 130350
rect 454058 130294 484598 130350
rect 484654 130294 484722 130350
rect 484778 130294 515318 130350
rect 515374 130294 515442 130350
rect 515498 130294 546038 130350
rect 546094 130294 546162 130350
rect 546218 130294 561250 130350
rect 561306 130294 561374 130350
rect 561430 130294 561498 130350
rect 561554 130294 561622 130350
rect 561678 130294 579250 130350
rect 579306 130294 579374 130350
rect 579430 130294 579498 130350
rect 579554 130294 579622 130350
rect 579678 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597980 130350
rect -1916 130226 597980 130294
rect -1916 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 3250 130226
rect 3306 130170 3374 130226
rect 3430 130170 3498 130226
rect 3554 130170 3622 130226
rect 3678 130170 21250 130226
rect 21306 130170 21374 130226
rect 21430 130170 21498 130226
rect 21554 130170 21622 130226
rect 21678 130170 39250 130226
rect 39306 130170 39374 130226
rect 39430 130170 39498 130226
rect 39554 130170 39622 130226
rect 39678 130170 54518 130226
rect 54574 130170 54642 130226
rect 54698 130170 57250 130226
rect 57306 130170 57374 130226
rect 57430 130170 57498 130226
rect 57554 130170 57622 130226
rect 57678 130170 75250 130226
rect 75306 130170 75374 130226
rect 75430 130170 75498 130226
rect 75554 130170 75622 130226
rect 75678 130170 85238 130226
rect 85294 130170 85362 130226
rect 85418 130170 93250 130226
rect 93306 130170 93374 130226
rect 93430 130170 93498 130226
rect 93554 130170 93622 130226
rect 93678 130170 111250 130226
rect 111306 130170 111374 130226
rect 111430 130170 111498 130226
rect 111554 130170 111622 130226
rect 111678 130170 115958 130226
rect 116014 130170 116082 130226
rect 116138 130170 146678 130226
rect 146734 130170 146802 130226
rect 146858 130170 177398 130226
rect 177454 130170 177522 130226
rect 177578 130170 208118 130226
rect 208174 130170 208242 130226
rect 208298 130170 238838 130226
rect 238894 130170 238962 130226
rect 239018 130170 269558 130226
rect 269614 130170 269682 130226
rect 269738 130170 300278 130226
rect 300334 130170 300402 130226
rect 300458 130170 330998 130226
rect 331054 130170 331122 130226
rect 331178 130170 361718 130226
rect 361774 130170 361842 130226
rect 361898 130170 392438 130226
rect 392494 130170 392562 130226
rect 392618 130170 423158 130226
rect 423214 130170 423282 130226
rect 423338 130170 453878 130226
rect 453934 130170 454002 130226
rect 454058 130170 484598 130226
rect 484654 130170 484722 130226
rect 484778 130170 515318 130226
rect 515374 130170 515442 130226
rect 515498 130170 546038 130226
rect 546094 130170 546162 130226
rect 546218 130170 561250 130226
rect 561306 130170 561374 130226
rect 561430 130170 561498 130226
rect 561554 130170 561622 130226
rect 561678 130170 579250 130226
rect 579306 130170 579374 130226
rect 579430 130170 579498 130226
rect 579554 130170 579622 130226
rect 579678 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597980 130226
rect -1916 130102 597980 130170
rect -1916 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 3250 130102
rect 3306 130046 3374 130102
rect 3430 130046 3498 130102
rect 3554 130046 3622 130102
rect 3678 130046 21250 130102
rect 21306 130046 21374 130102
rect 21430 130046 21498 130102
rect 21554 130046 21622 130102
rect 21678 130046 39250 130102
rect 39306 130046 39374 130102
rect 39430 130046 39498 130102
rect 39554 130046 39622 130102
rect 39678 130046 54518 130102
rect 54574 130046 54642 130102
rect 54698 130046 57250 130102
rect 57306 130046 57374 130102
rect 57430 130046 57498 130102
rect 57554 130046 57622 130102
rect 57678 130046 75250 130102
rect 75306 130046 75374 130102
rect 75430 130046 75498 130102
rect 75554 130046 75622 130102
rect 75678 130046 85238 130102
rect 85294 130046 85362 130102
rect 85418 130046 93250 130102
rect 93306 130046 93374 130102
rect 93430 130046 93498 130102
rect 93554 130046 93622 130102
rect 93678 130046 111250 130102
rect 111306 130046 111374 130102
rect 111430 130046 111498 130102
rect 111554 130046 111622 130102
rect 111678 130046 115958 130102
rect 116014 130046 116082 130102
rect 116138 130046 146678 130102
rect 146734 130046 146802 130102
rect 146858 130046 177398 130102
rect 177454 130046 177522 130102
rect 177578 130046 208118 130102
rect 208174 130046 208242 130102
rect 208298 130046 238838 130102
rect 238894 130046 238962 130102
rect 239018 130046 269558 130102
rect 269614 130046 269682 130102
rect 269738 130046 300278 130102
rect 300334 130046 300402 130102
rect 300458 130046 330998 130102
rect 331054 130046 331122 130102
rect 331178 130046 361718 130102
rect 361774 130046 361842 130102
rect 361898 130046 392438 130102
rect 392494 130046 392562 130102
rect 392618 130046 423158 130102
rect 423214 130046 423282 130102
rect 423338 130046 453878 130102
rect 453934 130046 454002 130102
rect 454058 130046 484598 130102
rect 484654 130046 484722 130102
rect 484778 130046 515318 130102
rect 515374 130046 515442 130102
rect 515498 130046 546038 130102
rect 546094 130046 546162 130102
rect 546218 130046 561250 130102
rect 561306 130046 561374 130102
rect 561430 130046 561498 130102
rect 561554 130046 561622 130102
rect 561678 130046 579250 130102
rect 579306 130046 579374 130102
rect 579430 130046 579498 130102
rect 579554 130046 579622 130102
rect 579678 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597980 130102
rect -1916 129978 597980 130046
rect -1916 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 3250 129978
rect 3306 129922 3374 129978
rect 3430 129922 3498 129978
rect 3554 129922 3622 129978
rect 3678 129922 21250 129978
rect 21306 129922 21374 129978
rect 21430 129922 21498 129978
rect 21554 129922 21622 129978
rect 21678 129922 39250 129978
rect 39306 129922 39374 129978
rect 39430 129922 39498 129978
rect 39554 129922 39622 129978
rect 39678 129922 54518 129978
rect 54574 129922 54642 129978
rect 54698 129922 57250 129978
rect 57306 129922 57374 129978
rect 57430 129922 57498 129978
rect 57554 129922 57622 129978
rect 57678 129922 75250 129978
rect 75306 129922 75374 129978
rect 75430 129922 75498 129978
rect 75554 129922 75622 129978
rect 75678 129922 85238 129978
rect 85294 129922 85362 129978
rect 85418 129922 93250 129978
rect 93306 129922 93374 129978
rect 93430 129922 93498 129978
rect 93554 129922 93622 129978
rect 93678 129922 111250 129978
rect 111306 129922 111374 129978
rect 111430 129922 111498 129978
rect 111554 129922 111622 129978
rect 111678 129922 115958 129978
rect 116014 129922 116082 129978
rect 116138 129922 146678 129978
rect 146734 129922 146802 129978
rect 146858 129922 177398 129978
rect 177454 129922 177522 129978
rect 177578 129922 208118 129978
rect 208174 129922 208242 129978
rect 208298 129922 238838 129978
rect 238894 129922 238962 129978
rect 239018 129922 269558 129978
rect 269614 129922 269682 129978
rect 269738 129922 300278 129978
rect 300334 129922 300402 129978
rect 300458 129922 330998 129978
rect 331054 129922 331122 129978
rect 331178 129922 361718 129978
rect 361774 129922 361842 129978
rect 361898 129922 392438 129978
rect 392494 129922 392562 129978
rect 392618 129922 423158 129978
rect 423214 129922 423282 129978
rect 423338 129922 453878 129978
rect 453934 129922 454002 129978
rect 454058 129922 484598 129978
rect 484654 129922 484722 129978
rect 484778 129922 515318 129978
rect 515374 129922 515442 129978
rect 515498 129922 546038 129978
rect 546094 129922 546162 129978
rect 546218 129922 561250 129978
rect 561306 129922 561374 129978
rect 561430 129922 561498 129978
rect 561554 129922 561622 129978
rect 561678 129922 579250 129978
rect 579306 129922 579374 129978
rect 579430 129922 579498 129978
rect 579554 129922 579622 129978
rect 579678 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597980 129978
rect -1916 129826 597980 129922
rect -1916 118350 597980 118446
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 6970 118350
rect 7026 118294 7094 118350
rect 7150 118294 7218 118350
rect 7274 118294 7342 118350
rect 7398 118294 24970 118350
rect 25026 118294 25094 118350
rect 25150 118294 25218 118350
rect 25274 118294 25342 118350
rect 25398 118294 42970 118350
rect 43026 118294 43094 118350
rect 43150 118294 43218 118350
rect 43274 118294 43342 118350
rect 43398 118294 60970 118350
rect 61026 118294 61094 118350
rect 61150 118294 61218 118350
rect 61274 118294 61342 118350
rect 61398 118294 69878 118350
rect 69934 118294 70002 118350
rect 70058 118294 78970 118350
rect 79026 118294 79094 118350
rect 79150 118294 79218 118350
rect 79274 118294 79342 118350
rect 79398 118294 96970 118350
rect 97026 118294 97094 118350
rect 97150 118294 97218 118350
rect 97274 118294 97342 118350
rect 97398 118294 100598 118350
rect 100654 118294 100722 118350
rect 100778 118294 131318 118350
rect 131374 118294 131442 118350
rect 131498 118294 162038 118350
rect 162094 118294 162162 118350
rect 162218 118294 192758 118350
rect 192814 118294 192882 118350
rect 192938 118294 223478 118350
rect 223534 118294 223602 118350
rect 223658 118294 254198 118350
rect 254254 118294 254322 118350
rect 254378 118294 284918 118350
rect 284974 118294 285042 118350
rect 285098 118294 315638 118350
rect 315694 118294 315762 118350
rect 315818 118294 346358 118350
rect 346414 118294 346482 118350
rect 346538 118294 377078 118350
rect 377134 118294 377202 118350
rect 377258 118294 407798 118350
rect 407854 118294 407922 118350
rect 407978 118294 438518 118350
rect 438574 118294 438642 118350
rect 438698 118294 469238 118350
rect 469294 118294 469362 118350
rect 469418 118294 499958 118350
rect 500014 118294 500082 118350
rect 500138 118294 530678 118350
rect 530734 118294 530802 118350
rect 530858 118294 564970 118350
rect 565026 118294 565094 118350
rect 565150 118294 565218 118350
rect 565274 118294 565342 118350
rect 565398 118294 582970 118350
rect 583026 118294 583094 118350
rect 583150 118294 583218 118350
rect 583274 118294 583342 118350
rect 583398 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect -1916 118226 597980 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 6970 118226
rect 7026 118170 7094 118226
rect 7150 118170 7218 118226
rect 7274 118170 7342 118226
rect 7398 118170 24970 118226
rect 25026 118170 25094 118226
rect 25150 118170 25218 118226
rect 25274 118170 25342 118226
rect 25398 118170 42970 118226
rect 43026 118170 43094 118226
rect 43150 118170 43218 118226
rect 43274 118170 43342 118226
rect 43398 118170 60970 118226
rect 61026 118170 61094 118226
rect 61150 118170 61218 118226
rect 61274 118170 61342 118226
rect 61398 118170 69878 118226
rect 69934 118170 70002 118226
rect 70058 118170 78970 118226
rect 79026 118170 79094 118226
rect 79150 118170 79218 118226
rect 79274 118170 79342 118226
rect 79398 118170 96970 118226
rect 97026 118170 97094 118226
rect 97150 118170 97218 118226
rect 97274 118170 97342 118226
rect 97398 118170 100598 118226
rect 100654 118170 100722 118226
rect 100778 118170 131318 118226
rect 131374 118170 131442 118226
rect 131498 118170 162038 118226
rect 162094 118170 162162 118226
rect 162218 118170 192758 118226
rect 192814 118170 192882 118226
rect 192938 118170 223478 118226
rect 223534 118170 223602 118226
rect 223658 118170 254198 118226
rect 254254 118170 254322 118226
rect 254378 118170 284918 118226
rect 284974 118170 285042 118226
rect 285098 118170 315638 118226
rect 315694 118170 315762 118226
rect 315818 118170 346358 118226
rect 346414 118170 346482 118226
rect 346538 118170 377078 118226
rect 377134 118170 377202 118226
rect 377258 118170 407798 118226
rect 407854 118170 407922 118226
rect 407978 118170 438518 118226
rect 438574 118170 438642 118226
rect 438698 118170 469238 118226
rect 469294 118170 469362 118226
rect 469418 118170 499958 118226
rect 500014 118170 500082 118226
rect 500138 118170 530678 118226
rect 530734 118170 530802 118226
rect 530858 118170 564970 118226
rect 565026 118170 565094 118226
rect 565150 118170 565218 118226
rect 565274 118170 565342 118226
rect 565398 118170 582970 118226
rect 583026 118170 583094 118226
rect 583150 118170 583218 118226
rect 583274 118170 583342 118226
rect 583398 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect -1916 118102 597980 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 6970 118102
rect 7026 118046 7094 118102
rect 7150 118046 7218 118102
rect 7274 118046 7342 118102
rect 7398 118046 24970 118102
rect 25026 118046 25094 118102
rect 25150 118046 25218 118102
rect 25274 118046 25342 118102
rect 25398 118046 42970 118102
rect 43026 118046 43094 118102
rect 43150 118046 43218 118102
rect 43274 118046 43342 118102
rect 43398 118046 60970 118102
rect 61026 118046 61094 118102
rect 61150 118046 61218 118102
rect 61274 118046 61342 118102
rect 61398 118046 69878 118102
rect 69934 118046 70002 118102
rect 70058 118046 78970 118102
rect 79026 118046 79094 118102
rect 79150 118046 79218 118102
rect 79274 118046 79342 118102
rect 79398 118046 96970 118102
rect 97026 118046 97094 118102
rect 97150 118046 97218 118102
rect 97274 118046 97342 118102
rect 97398 118046 100598 118102
rect 100654 118046 100722 118102
rect 100778 118046 131318 118102
rect 131374 118046 131442 118102
rect 131498 118046 162038 118102
rect 162094 118046 162162 118102
rect 162218 118046 192758 118102
rect 192814 118046 192882 118102
rect 192938 118046 223478 118102
rect 223534 118046 223602 118102
rect 223658 118046 254198 118102
rect 254254 118046 254322 118102
rect 254378 118046 284918 118102
rect 284974 118046 285042 118102
rect 285098 118046 315638 118102
rect 315694 118046 315762 118102
rect 315818 118046 346358 118102
rect 346414 118046 346482 118102
rect 346538 118046 377078 118102
rect 377134 118046 377202 118102
rect 377258 118046 407798 118102
rect 407854 118046 407922 118102
rect 407978 118046 438518 118102
rect 438574 118046 438642 118102
rect 438698 118046 469238 118102
rect 469294 118046 469362 118102
rect 469418 118046 499958 118102
rect 500014 118046 500082 118102
rect 500138 118046 530678 118102
rect 530734 118046 530802 118102
rect 530858 118046 564970 118102
rect 565026 118046 565094 118102
rect 565150 118046 565218 118102
rect 565274 118046 565342 118102
rect 565398 118046 582970 118102
rect 583026 118046 583094 118102
rect 583150 118046 583218 118102
rect 583274 118046 583342 118102
rect 583398 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect -1916 117978 597980 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 6970 117978
rect 7026 117922 7094 117978
rect 7150 117922 7218 117978
rect 7274 117922 7342 117978
rect 7398 117922 24970 117978
rect 25026 117922 25094 117978
rect 25150 117922 25218 117978
rect 25274 117922 25342 117978
rect 25398 117922 42970 117978
rect 43026 117922 43094 117978
rect 43150 117922 43218 117978
rect 43274 117922 43342 117978
rect 43398 117922 60970 117978
rect 61026 117922 61094 117978
rect 61150 117922 61218 117978
rect 61274 117922 61342 117978
rect 61398 117922 69878 117978
rect 69934 117922 70002 117978
rect 70058 117922 78970 117978
rect 79026 117922 79094 117978
rect 79150 117922 79218 117978
rect 79274 117922 79342 117978
rect 79398 117922 96970 117978
rect 97026 117922 97094 117978
rect 97150 117922 97218 117978
rect 97274 117922 97342 117978
rect 97398 117922 100598 117978
rect 100654 117922 100722 117978
rect 100778 117922 131318 117978
rect 131374 117922 131442 117978
rect 131498 117922 162038 117978
rect 162094 117922 162162 117978
rect 162218 117922 192758 117978
rect 192814 117922 192882 117978
rect 192938 117922 223478 117978
rect 223534 117922 223602 117978
rect 223658 117922 254198 117978
rect 254254 117922 254322 117978
rect 254378 117922 284918 117978
rect 284974 117922 285042 117978
rect 285098 117922 315638 117978
rect 315694 117922 315762 117978
rect 315818 117922 346358 117978
rect 346414 117922 346482 117978
rect 346538 117922 377078 117978
rect 377134 117922 377202 117978
rect 377258 117922 407798 117978
rect 407854 117922 407922 117978
rect 407978 117922 438518 117978
rect 438574 117922 438642 117978
rect 438698 117922 469238 117978
rect 469294 117922 469362 117978
rect 469418 117922 499958 117978
rect 500014 117922 500082 117978
rect 500138 117922 530678 117978
rect 530734 117922 530802 117978
rect 530858 117922 564970 117978
rect 565026 117922 565094 117978
rect 565150 117922 565218 117978
rect 565274 117922 565342 117978
rect 565398 117922 582970 117978
rect 583026 117922 583094 117978
rect 583150 117922 583218 117978
rect 583274 117922 583342 117978
rect 583398 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect -1916 117826 597980 117922
rect -1916 112350 597980 112446
rect -1916 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 3250 112350
rect 3306 112294 3374 112350
rect 3430 112294 3498 112350
rect 3554 112294 3622 112350
rect 3678 112294 21250 112350
rect 21306 112294 21374 112350
rect 21430 112294 21498 112350
rect 21554 112294 21622 112350
rect 21678 112294 39250 112350
rect 39306 112294 39374 112350
rect 39430 112294 39498 112350
rect 39554 112294 39622 112350
rect 39678 112294 54518 112350
rect 54574 112294 54642 112350
rect 54698 112294 57250 112350
rect 57306 112294 57374 112350
rect 57430 112294 57498 112350
rect 57554 112294 57622 112350
rect 57678 112294 75250 112350
rect 75306 112294 75374 112350
rect 75430 112294 75498 112350
rect 75554 112294 75622 112350
rect 75678 112294 85238 112350
rect 85294 112294 85362 112350
rect 85418 112294 93250 112350
rect 93306 112294 93374 112350
rect 93430 112294 93498 112350
rect 93554 112294 93622 112350
rect 93678 112294 111250 112350
rect 111306 112294 111374 112350
rect 111430 112294 111498 112350
rect 111554 112294 111622 112350
rect 111678 112294 115958 112350
rect 116014 112294 116082 112350
rect 116138 112294 146678 112350
rect 146734 112294 146802 112350
rect 146858 112294 177398 112350
rect 177454 112294 177522 112350
rect 177578 112294 208118 112350
rect 208174 112294 208242 112350
rect 208298 112294 238838 112350
rect 238894 112294 238962 112350
rect 239018 112294 269558 112350
rect 269614 112294 269682 112350
rect 269738 112294 300278 112350
rect 300334 112294 300402 112350
rect 300458 112294 330998 112350
rect 331054 112294 331122 112350
rect 331178 112294 361718 112350
rect 361774 112294 361842 112350
rect 361898 112294 392438 112350
rect 392494 112294 392562 112350
rect 392618 112294 423158 112350
rect 423214 112294 423282 112350
rect 423338 112294 453878 112350
rect 453934 112294 454002 112350
rect 454058 112294 484598 112350
rect 484654 112294 484722 112350
rect 484778 112294 515318 112350
rect 515374 112294 515442 112350
rect 515498 112294 546038 112350
rect 546094 112294 546162 112350
rect 546218 112294 561250 112350
rect 561306 112294 561374 112350
rect 561430 112294 561498 112350
rect 561554 112294 561622 112350
rect 561678 112294 579250 112350
rect 579306 112294 579374 112350
rect 579430 112294 579498 112350
rect 579554 112294 579622 112350
rect 579678 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597980 112350
rect -1916 112226 597980 112294
rect -1916 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 3250 112226
rect 3306 112170 3374 112226
rect 3430 112170 3498 112226
rect 3554 112170 3622 112226
rect 3678 112170 21250 112226
rect 21306 112170 21374 112226
rect 21430 112170 21498 112226
rect 21554 112170 21622 112226
rect 21678 112170 39250 112226
rect 39306 112170 39374 112226
rect 39430 112170 39498 112226
rect 39554 112170 39622 112226
rect 39678 112170 54518 112226
rect 54574 112170 54642 112226
rect 54698 112170 57250 112226
rect 57306 112170 57374 112226
rect 57430 112170 57498 112226
rect 57554 112170 57622 112226
rect 57678 112170 75250 112226
rect 75306 112170 75374 112226
rect 75430 112170 75498 112226
rect 75554 112170 75622 112226
rect 75678 112170 85238 112226
rect 85294 112170 85362 112226
rect 85418 112170 93250 112226
rect 93306 112170 93374 112226
rect 93430 112170 93498 112226
rect 93554 112170 93622 112226
rect 93678 112170 111250 112226
rect 111306 112170 111374 112226
rect 111430 112170 111498 112226
rect 111554 112170 111622 112226
rect 111678 112170 115958 112226
rect 116014 112170 116082 112226
rect 116138 112170 146678 112226
rect 146734 112170 146802 112226
rect 146858 112170 177398 112226
rect 177454 112170 177522 112226
rect 177578 112170 208118 112226
rect 208174 112170 208242 112226
rect 208298 112170 238838 112226
rect 238894 112170 238962 112226
rect 239018 112170 269558 112226
rect 269614 112170 269682 112226
rect 269738 112170 300278 112226
rect 300334 112170 300402 112226
rect 300458 112170 330998 112226
rect 331054 112170 331122 112226
rect 331178 112170 361718 112226
rect 361774 112170 361842 112226
rect 361898 112170 392438 112226
rect 392494 112170 392562 112226
rect 392618 112170 423158 112226
rect 423214 112170 423282 112226
rect 423338 112170 453878 112226
rect 453934 112170 454002 112226
rect 454058 112170 484598 112226
rect 484654 112170 484722 112226
rect 484778 112170 515318 112226
rect 515374 112170 515442 112226
rect 515498 112170 546038 112226
rect 546094 112170 546162 112226
rect 546218 112170 561250 112226
rect 561306 112170 561374 112226
rect 561430 112170 561498 112226
rect 561554 112170 561622 112226
rect 561678 112170 579250 112226
rect 579306 112170 579374 112226
rect 579430 112170 579498 112226
rect 579554 112170 579622 112226
rect 579678 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597980 112226
rect -1916 112102 597980 112170
rect -1916 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 3250 112102
rect 3306 112046 3374 112102
rect 3430 112046 3498 112102
rect 3554 112046 3622 112102
rect 3678 112046 21250 112102
rect 21306 112046 21374 112102
rect 21430 112046 21498 112102
rect 21554 112046 21622 112102
rect 21678 112046 39250 112102
rect 39306 112046 39374 112102
rect 39430 112046 39498 112102
rect 39554 112046 39622 112102
rect 39678 112046 54518 112102
rect 54574 112046 54642 112102
rect 54698 112046 57250 112102
rect 57306 112046 57374 112102
rect 57430 112046 57498 112102
rect 57554 112046 57622 112102
rect 57678 112046 75250 112102
rect 75306 112046 75374 112102
rect 75430 112046 75498 112102
rect 75554 112046 75622 112102
rect 75678 112046 85238 112102
rect 85294 112046 85362 112102
rect 85418 112046 93250 112102
rect 93306 112046 93374 112102
rect 93430 112046 93498 112102
rect 93554 112046 93622 112102
rect 93678 112046 111250 112102
rect 111306 112046 111374 112102
rect 111430 112046 111498 112102
rect 111554 112046 111622 112102
rect 111678 112046 115958 112102
rect 116014 112046 116082 112102
rect 116138 112046 146678 112102
rect 146734 112046 146802 112102
rect 146858 112046 177398 112102
rect 177454 112046 177522 112102
rect 177578 112046 208118 112102
rect 208174 112046 208242 112102
rect 208298 112046 238838 112102
rect 238894 112046 238962 112102
rect 239018 112046 269558 112102
rect 269614 112046 269682 112102
rect 269738 112046 300278 112102
rect 300334 112046 300402 112102
rect 300458 112046 330998 112102
rect 331054 112046 331122 112102
rect 331178 112046 361718 112102
rect 361774 112046 361842 112102
rect 361898 112046 392438 112102
rect 392494 112046 392562 112102
rect 392618 112046 423158 112102
rect 423214 112046 423282 112102
rect 423338 112046 453878 112102
rect 453934 112046 454002 112102
rect 454058 112046 484598 112102
rect 484654 112046 484722 112102
rect 484778 112046 515318 112102
rect 515374 112046 515442 112102
rect 515498 112046 546038 112102
rect 546094 112046 546162 112102
rect 546218 112046 561250 112102
rect 561306 112046 561374 112102
rect 561430 112046 561498 112102
rect 561554 112046 561622 112102
rect 561678 112046 579250 112102
rect 579306 112046 579374 112102
rect 579430 112046 579498 112102
rect 579554 112046 579622 112102
rect 579678 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597980 112102
rect -1916 111978 597980 112046
rect -1916 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 3250 111978
rect 3306 111922 3374 111978
rect 3430 111922 3498 111978
rect 3554 111922 3622 111978
rect 3678 111922 21250 111978
rect 21306 111922 21374 111978
rect 21430 111922 21498 111978
rect 21554 111922 21622 111978
rect 21678 111922 39250 111978
rect 39306 111922 39374 111978
rect 39430 111922 39498 111978
rect 39554 111922 39622 111978
rect 39678 111922 54518 111978
rect 54574 111922 54642 111978
rect 54698 111922 57250 111978
rect 57306 111922 57374 111978
rect 57430 111922 57498 111978
rect 57554 111922 57622 111978
rect 57678 111922 75250 111978
rect 75306 111922 75374 111978
rect 75430 111922 75498 111978
rect 75554 111922 75622 111978
rect 75678 111922 85238 111978
rect 85294 111922 85362 111978
rect 85418 111922 93250 111978
rect 93306 111922 93374 111978
rect 93430 111922 93498 111978
rect 93554 111922 93622 111978
rect 93678 111922 111250 111978
rect 111306 111922 111374 111978
rect 111430 111922 111498 111978
rect 111554 111922 111622 111978
rect 111678 111922 115958 111978
rect 116014 111922 116082 111978
rect 116138 111922 146678 111978
rect 146734 111922 146802 111978
rect 146858 111922 177398 111978
rect 177454 111922 177522 111978
rect 177578 111922 208118 111978
rect 208174 111922 208242 111978
rect 208298 111922 238838 111978
rect 238894 111922 238962 111978
rect 239018 111922 269558 111978
rect 269614 111922 269682 111978
rect 269738 111922 300278 111978
rect 300334 111922 300402 111978
rect 300458 111922 330998 111978
rect 331054 111922 331122 111978
rect 331178 111922 361718 111978
rect 361774 111922 361842 111978
rect 361898 111922 392438 111978
rect 392494 111922 392562 111978
rect 392618 111922 423158 111978
rect 423214 111922 423282 111978
rect 423338 111922 453878 111978
rect 453934 111922 454002 111978
rect 454058 111922 484598 111978
rect 484654 111922 484722 111978
rect 484778 111922 515318 111978
rect 515374 111922 515442 111978
rect 515498 111922 546038 111978
rect 546094 111922 546162 111978
rect 546218 111922 561250 111978
rect 561306 111922 561374 111978
rect 561430 111922 561498 111978
rect 561554 111922 561622 111978
rect 561678 111922 579250 111978
rect 579306 111922 579374 111978
rect 579430 111922 579498 111978
rect 579554 111922 579622 111978
rect 579678 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597980 111978
rect -1916 111826 597980 111922
rect -1916 100350 597980 100446
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 6970 100350
rect 7026 100294 7094 100350
rect 7150 100294 7218 100350
rect 7274 100294 7342 100350
rect 7398 100294 24970 100350
rect 25026 100294 25094 100350
rect 25150 100294 25218 100350
rect 25274 100294 25342 100350
rect 25398 100294 42970 100350
rect 43026 100294 43094 100350
rect 43150 100294 43218 100350
rect 43274 100294 43342 100350
rect 43398 100294 60970 100350
rect 61026 100294 61094 100350
rect 61150 100294 61218 100350
rect 61274 100294 61342 100350
rect 61398 100294 69878 100350
rect 69934 100294 70002 100350
rect 70058 100294 78970 100350
rect 79026 100294 79094 100350
rect 79150 100294 79218 100350
rect 79274 100294 79342 100350
rect 79398 100294 96970 100350
rect 97026 100294 97094 100350
rect 97150 100294 97218 100350
rect 97274 100294 97342 100350
rect 97398 100294 100598 100350
rect 100654 100294 100722 100350
rect 100778 100294 131318 100350
rect 131374 100294 131442 100350
rect 131498 100294 162038 100350
rect 162094 100294 162162 100350
rect 162218 100294 192758 100350
rect 192814 100294 192882 100350
rect 192938 100294 223478 100350
rect 223534 100294 223602 100350
rect 223658 100294 254198 100350
rect 254254 100294 254322 100350
rect 254378 100294 284918 100350
rect 284974 100294 285042 100350
rect 285098 100294 315638 100350
rect 315694 100294 315762 100350
rect 315818 100294 346358 100350
rect 346414 100294 346482 100350
rect 346538 100294 377078 100350
rect 377134 100294 377202 100350
rect 377258 100294 407798 100350
rect 407854 100294 407922 100350
rect 407978 100294 438518 100350
rect 438574 100294 438642 100350
rect 438698 100294 469238 100350
rect 469294 100294 469362 100350
rect 469418 100294 499958 100350
rect 500014 100294 500082 100350
rect 500138 100294 530678 100350
rect 530734 100294 530802 100350
rect 530858 100294 564970 100350
rect 565026 100294 565094 100350
rect 565150 100294 565218 100350
rect 565274 100294 565342 100350
rect 565398 100294 582970 100350
rect 583026 100294 583094 100350
rect 583150 100294 583218 100350
rect 583274 100294 583342 100350
rect 583398 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect -1916 100226 597980 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 6970 100226
rect 7026 100170 7094 100226
rect 7150 100170 7218 100226
rect 7274 100170 7342 100226
rect 7398 100170 24970 100226
rect 25026 100170 25094 100226
rect 25150 100170 25218 100226
rect 25274 100170 25342 100226
rect 25398 100170 42970 100226
rect 43026 100170 43094 100226
rect 43150 100170 43218 100226
rect 43274 100170 43342 100226
rect 43398 100170 60970 100226
rect 61026 100170 61094 100226
rect 61150 100170 61218 100226
rect 61274 100170 61342 100226
rect 61398 100170 69878 100226
rect 69934 100170 70002 100226
rect 70058 100170 78970 100226
rect 79026 100170 79094 100226
rect 79150 100170 79218 100226
rect 79274 100170 79342 100226
rect 79398 100170 96970 100226
rect 97026 100170 97094 100226
rect 97150 100170 97218 100226
rect 97274 100170 97342 100226
rect 97398 100170 100598 100226
rect 100654 100170 100722 100226
rect 100778 100170 131318 100226
rect 131374 100170 131442 100226
rect 131498 100170 162038 100226
rect 162094 100170 162162 100226
rect 162218 100170 192758 100226
rect 192814 100170 192882 100226
rect 192938 100170 223478 100226
rect 223534 100170 223602 100226
rect 223658 100170 254198 100226
rect 254254 100170 254322 100226
rect 254378 100170 284918 100226
rect 284974 100170 285042 100226
rect 285098 100170 315638 100226
rect 315694 100170 315762 100226
rect 315818 100170 346358 100226
rect 346414 100170 346482 100226
rect 346538 100170 377078 100226
rect 377134 100170 377202 100226
rect 377258 100170 407798 100226
rect 407854 100170 407922 100226
rect 407978 100170 438518 100226
rect 438574 100170 438642 100226
rect 438698 100170 469238 100226
rect 469294 100170 469362 100226
rect 469418 100170 499958 100226
rect 500014 100170 500082 100226
rect 500138 100170 530678 100226
rect 530734 100170 530802 100226
rect 530858 100170 564970 100226
rect 565026 100170 565094 100226
rect 565150 100170 565218 100226
rect 565274 100170 565342 100226
rect 565398 100170 582970 100226
rect 583026 100170 583094 100226
rect 583150 100170 583218 100226
rect 583274 100170 583342 100226
rect 583398 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect -1916 100102 597980 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 6970 100102
rect 7026 100046 7094 100102
rect 7150 100046 7218 100102
rect 7274 100046 7342 100102
rect 7398 100046 24970 100102
rect 25026 100046 25094 100102
rect 25150 100046 25218 100102
rect 25274 100046 25342 100102
rect 25398 100046 42970 100102
rect 43026 100046 43094 100102
rect 43150 100046 43218 100102
rect 43274 100046 43342 100102
rect 43398 100046 60970 100102
rect 61026 100046 61094 100102
rect 61150 100046 61218 100102
rect 61274 100046 61342 100102
rect 61398 100046 69878 100102
rect 69934 100046 70002 100102
rect 70058 100046 78970 100102
rect 79026 100046 79094 100102
rect 79150 100046 79218 100102
rect 79274 100046 79342 100102
rect 79398 100046 96970 100102
rect 97026 100046 97094 100102
rect 97150 100046 97218 100102
rect 97274 100046 97342 100102
rect 97398 100046 100598 100102
rect 100654 100046 100722 100102
rect 100778 100046 131318 100102
rect 131374 100046 131442 100102
rect 131498 100046 162038 100102
rect 162094 100046 162162 100102
rect 162218 100046 192758 100102
rect 192814 100046 192882 100102
rect 192938 100046 223478 100102
rect 223534 100046 223602 100102
rect 223658 100046 254198 100102
rect 254254 100046 254322 100102
rect 254378 100046 284918 100102
rect 284974 100046 285042 100102
rect 285098 100046 315638 100102
rect 315694 100046 315762 100102
rect 315818 100046 346358 100102
rect 346414 100046 346482 100102
rect 346538 100046 377078 100102
rect 377134 100046 377202 100102
rect 377258 100046 407798 100102
rect 407854 100046 407922 100102
rect 407978 100046 438518 100102
rect 438574 100046 438642 100102
rect 438698 100046 469238 100102
rect 469294 100046 469362 100102
rect 469418 100046 499958 100102
rect 500014 100046 500082 100102
rect 500138 100046 530678 100102
rect 530734 100046 530802 100102
rect 530858 100046 564970 100102
rect 565026 100046 565094 100102
rect 565150 100046 565218 100102
rect 565274 100046 565342 100102
rect 565398 100046 582970 100102
rect 583026 100046 583094 100102
rect 583150 100046 583218 100102
rect 583274 100046 583342 100102
rect 583398 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect -1916 99978 597980 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 6970 99978
rect 7026 99922 7094 99978
rect 7150 99922 7218 99978
rect 7274 99922 7342 99978
rect 7398 99922 24970 99978
rect 25026 99922 25094 99978
rect 25150 99922 25218 99978
rect 25274 99922 25342 99978
rect 25398 99922 42970 99978
rect 43026 99922 43094 99978
rect 43150 99922 43218 99978
rect 43274 99922 43342 99978
rect 43398 99922 60970 99978
rect 61026 99922 61094 99978
rect 61150 99922 61218 99978
rect 61274 99922 61342 99978
rect 61398 99922 69878 99978
rect 69934 99922 70002 99978
rect 70058 99922 78970 99978
rect 79026 99922 79094 99978
rect 79150 99922 79218 99978
rect 79274 99922 79342 99978
rect 79398 99922 96970 99978
rect 97026 99922 97094 99978
rect 97150 99922 97218 99978
rect 97274 99922 97342 99978
rect 97398 99922 100598 99978
rect 100654 99922 100722 99978
rect 100778 99922 131318 99978
rect 131374 99922 131442 99978
rect 131498 99922 162038 99978
rect 162094 99922 162162 99978
rect 162218 99922 192758 99978
rect 192814 99922 192882 99978
rect 192938 99922 223478 99978
rect 223534 99922 223602 99978
rect 223658 99922 254198 99978
rect 254254 99922 254322 99978
rect 254378 99922 284918 99978
rect 284974 99922 285042 99978
rect 285098 99922 315638 99978
rect 315694 99922 315762 99978
rect 315818 99922 346358 99978
rect 346414 99922 346482 99978
rect 346538 99922 377078 99978
rect 377134 99922 377202 99978
rect 377258 99922 407798 99978
rect 407854 99922 407922 99978
rect 407978 99922 438518 99978
rect 438574 99922 438642 99978
rect 438698 99922 469238 99978
rect 469294 99922 469362 99978
rect 469418 99922 499958 99978
rect 500014 99922 500082 99978
rect 500138 99922 530678 99978
rect 530734 99922 530802 99978
rect 530858 99922 564970 99978
rect 565026 99922 565094 99978
rect 565150 99922 565218 99978
rect 565274 99922 565342 99978
rect 565398 99922 582970 99978
rect 583026 99922 583094 99978
rect 583150 99922 583218 99978
rect 583274 99922 583342 99978
rect 583398 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect -1916 99826 597980 99922
rect -1916 94350 597980 94446
rect -1916 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 3250 94350
rect 3306 94294 3374 94350
rect 3430 94294 3498 94350
rect 3554 94294 3622 94350
rect 3678 94294 21250 94350
rect 21306 94294 21374 94350
rect 21430 94294 21498 94350
rect 21554 94294 21622 94350
rect 21678 94294 39250 94350
rect 39306 94294 39374 94350
rect 39430 94294 39498 94350
rect 39554 94294 39622 94350
rect 39678 94294 54518 94350
rect 54574 94294 54642 94350
rect 54698 94294 57250 94350
rect 57306 94294 57374 94350
rect 57430 94294 57498 94350
rect 57554 94294 57622 94350
rect 57678 94294 75250 94350
rect 75306 94294 75374 94350
rect 75430 94294 75498 94350
rect 75554 94294 75622 94350
rect 75678 94294 85238 94350
rect 85294 94294 85362 94350
rect 85418 94294 93250 94350
rect 93306 94294 93374 94350
rect 93430 94294 93498 94350
rect 93554 94294 93622 94350
rect 93678 94294 111250 94350
rect 111306 94294 111374 94350
rect 111430 94294 111498 94350
rect 111554 94294 111622 94350
rect 111678 94294 115958 94350
rect 116014 94294 116082 94350
rect 116138 94294 146678 94350
rect 146734 94294 146802 94350
rect 146858 94294 177398 94350
rect 177454 94294 177522 94350
rect 177578 94294 208118 94350
rect 208174 94294 208242 94350
rect 208298 94294 238838 94350
rect 238894 94294 238962 94350
rect 239018 94294 269558 94350
rect 269614 94294 269682 94350
rect 269738 94294 300278 94350
rect 300334 94294 300402 94350
rect 300458 94294 330998 94350
rect 331054 94294 331122 94350
rect 331178 94294 361718 94350
rect 361774 94294 361842 94350
rect 361898 94294 392438 94350
rect 392494 94294 392562 94350
rect 392618 94294 423158 94350
rect 423214 94294 423282 94350
rect 423338 94294 453878 94350
rect 453934 94294 454002 94350
rect 454058 94294 484598 94350
rect 484654 94294 484722 94350
rect 484778 94294 515318 94350
rect 515374 94294 515442 94350
rect 515498 94294 546038 94350
rect 546094 94294 546162 94350
rect 546218 94294 561250 94350
rect 561306 94294 561374 94350
rect 561430 94294 561498 94350
rect 561554 94294 561622 94350
rect 561678 94294 579250 94350
rect 579306 94294 579374 94350
rect 579430 94294 579498 94350
rect 579554 94294 579622 94350
rect 579678 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597980 94350
rect -1916 94226 597980 94294
rect -1916 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 3250 94226
rect 3306 94170 3374 94226
rect 3430 94170 3498 94226
rect 3554 94170 3622 94226
rect 3678 94170 21250 94226
rect 21306 94170 21374 94226
rect 21430 94170 21498 94226
rect 21554 94170 21622 94226
rect 21678 94170 39250 94226
rect 39306 94170 39374 94226
rect 39430 94170 39498 94226
rect 39554 94170 39622 94226
rect 39678 94170 54518 94226
rect 54574 94170 54642 94226
rect 54698 94170 57250 94226
rect 57306 94170 57374 94226
rect 57430 94170 57498 94226
rect 57554 94170 57622 94226
rect 57678 94170 75250 94226
rect 75306 94170 75374 94226
rect 75430 94170 75498 94226
rect 75554 94170 75622 94226
rect 75678 94170 85238 94226
rect 85294 94170 85362 94226
rect 85418 94170 93250 94226
rect 93306 94170 93374 94226
rect 93430 94170 93498 94226
rect 93554 94170 93622 94226
rect 93678 94170 111250 94226
rect 111306 94170 111374 94226
rect 111430 94170 111498 94226
rect 111554 94170 111622 94226
rect 111678 94170 115958 94226
rect 116014 94170 116082 94226
rect 116138 94170 146678 94226
rect 146734 94170 146802 94226
rect 146858 94170 177398 94226
rect 177454 94170 177522 94226
rect 177578 94170 208118 94226
rect 208174 94170 208242 94226
rect 208298 94170 238838 94226
rect 238894 94170 238962 94226
rect 239018 94170 269558 94226
rect 269614 94170 269682 94226
rect 269738 94170 300278 94226
rect 300334 94170 300402 94226
rect 300458 94170 330998 94226
rect 331054 94170 331122 94226
rect 331178 94170 361718 94226
rect 361774 94170 361842 94226
rect 361898 94170 392438 94226
rect 392494 94170 392562 94226
rect 392618 94170 423158 94226
rect 423214 94170 423282 94226
rect 423338 94170 453878 94226
rect 453934 94170 454002 94226
rect 454058 94170 484598 94226
rect 484654 94170 484722 94226
rect 484778 94170 515318 94226
rect 515374 94170 515442 94226
rect 515498 94170 546038 94226
rect 546094 94170 546162 94226
rect 546218 94170 561250 94226
rect 561306 94170 561374 94226
rect 561430 94170 561498 94226
rect 561554 94170 561622 94226
rect 561678 94170 579250 94226
rect 579306 94170 579374 94226
rect 579430 94170 579498 94226
rect 579554 94170 579622 94226
rect 579678 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597980 94226
rect -1916 94102 597980 94170
rect -1916 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 3250 94102
rect 3306 94046 3374 94102
rect 3430 94046 3498 94102
rect 3554 94046 3622 94102
rect 3678 94046 21250 94102
rect 21306 94046 21374 94102
rect 21430 94046 21498 94102
rect 21554 94046 21622 94102
rect 21678 94046 39250 94102
rect 39306 94046 39374 94102
rect 39430 94046 39498 94102
rect 39554 94046 39622 94102
rect 39678 94046 54518 94102
rect 54574 94046 54642 94102
rect 54698 94046 57250 94102
rect 57306 94046 57374 94102
rect 57430 94046 57498 94102
rect 57554 94046 57622 94102
rect 57678 94046 75250 94102
rect 75306 94046 75374 94102
rect 75430 94046 75498 94102
rect 75554 94046 75622 94102
rect 75678 94046 85238 94102
rect 85294 94046 85362 94102
rect 85418 94046 93250 94102
rect 93306 94046 93374 94102
rect 93430 94046 93498 94102
rect 93554 94046 93622 94102
rect 93678 94046 111250 94102
rect 111306 94046 111374 94102
rect 111430 94046 111498 94102
rect 111554 94046 111622 94102
rect 111678 94046 115958 94102
rect 116014 94046 116082 94102
rect 116138 94046 146678 94102
rect 146734 94046 146802 94102
rect 146858 94046 177398 94102
rect 177454 94046 177522 94102
rect 177578 94046 208118 94102
rect 208174 94046 208242 94102
rect 208298 94046 238838 94102
rect 238894 94046 238962 94102
rect 239018 94046 269558 94102
rect 269614 94046 269682 94102
rect 269738 94046 300278 94102
rect 300334 94046 300402 94102
rect 300458 94046 330998 94102
rect 331054 94046 331122 94102
rect 331178 94046 361718 94102
rect 361774 94046 361842 94102
rect 361898 94046 392438 94102
rect 392494 94046 392562 94102
rect 392618 94046 423158 94102
rect 423214 94046 423282 94102
rect 423338 94046 453878 94102
rect 453934 94046 454002 94102
rect 454058 94046 484598 94102
rect 484654 94046 484722 94102
rect 484778 94046 515318 94102
rect 515374 94046 515442 94102
rect 515498 94046 546038 94102
rect 546094 94046 546162 94102
rect 546218 94046 561250 94102
rect 561306 94046 561374 94102
rect 561430 94046 561498 94102
rect 561554 94046 561622 94102
rect 561678 94046 579250 94102
rect 579306 94046 579374 94102
rect 579430 94046 579498 94102
rect 579554 94046 579622 94102
rect 579678 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597980 94102
rect -1916 93978 597980 94046
rect -1916 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 3250 93978
rect 3306 93922 3374 93978
rect 3430 93922 3498 93978
rect 3554 93922 3622 93978
rect 3678 93922 21250 93978
rect 21306 93922 21374 93978
rect 21430 93922 21498 93978
rect 21554 93922 21622 93978
rect 21678 93922 39250 93978
rect 39306 93922 39374 93978
rect 39430 93922 39498 93978
rect 39554 93922 39622 93978
rect 39678 93922 54518 93978
rect 54574 93922 54642 93978
rect 54698 93922 57250 93978
rect 57306 93922 57374 93978
rect 57430 93922 57498 93978
rect 57554 93922 57622 93978
rect 57678 93922 75250 93978
rect 75306 93922 75374 93978
rect 75430 93922 75498 93978
rect 75554 93922 75622 93978
rect 75678 93922 85238 93978
rect 85294 93922 85362 93978
rect 85418 93922 93250 93978
rect 93306 93922 93374 93978
rect 93430 93922 93498 93978
rect 93554 93922 93622 93978
rect 93678 93922 111250 93978
rect 111306 93922 111374 93978
rect 111430 93922 111498 93978
rect 111554 93922 111622 93978
rect 111678 93922 115958 93978
rect 116014 93922 116082 93978
rect 116138 93922 146678 93978
rect 146734 93922 146802 93978
rect 146858 93922 177398 93978
rect 177454 93922 177522 93978
rect 177578 93922 208118 93978
rect 208174 93922 208242 93978
rect 208298 93922 238838 93978
rect 238894 93922 238962 93978
rect 239018 93922 269558 93978
rect 269614 93922 269682 93978
rect 269738 93922 300278 93978
rect 300334 93922 300402 93978
rect 300458 93922 330998 93978
rect 331054 93922 331122 93978
rect 331178 93922 361718 93978
rect 361774 93922 361842 93978
rect 361898 93922 392438 93978
rect 392494 93922 392562 93978
rect 392618 93922 423158 93978
rect 423214 93922 423282 93978
rect 423338 93922 453878 93978
rect 453934 93922 454002 93978
rect 454058 93922 484598 93978
rect 484654 93922 484722 93978
rect 484778 93922 515318 93978
rect 515374 93922 515442 93978
rect 515498 93922 546038 93978
rect 546094 93922 546162 93978
rect 546218 93922 561250 93978
rect 561306 93922 561374 93978
rect 561430 93922 561498 93978
rect 561554 93922 561622 93978
rect 561678 93922 579250 93978
rect 579306 93922 579374 93978
rect 579430 93922 579498 93978
rect 579554 93922 579622 93978
rect 579678 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597980 93978
rect -1916 93826 597980 93922
rect -1916 82350 597980 82446
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 6970 82350
rect 7026 82294 7094 82350
rect 7150 82294 7218 82350
rect 7274 82294 7342 82350
rect 7398 82294 24970 82350
rect 25026 82294 25094 82350
rect 25150 82294 25218 82350
rect 25274 82294 25342 82350
rect 25398 82294 42970 82350
rect 43026 82294 43094 82350
rect 43150 82294 43218 82350
rect 43274 82294 43342 82350
rect 43398 82294 60970 82350
rect 61026 82294 61094 82350
rect 61150 82294 61218 82350
rect 61274 82294 61342 82350
rect 61398 82294 69878 82350
rect 69934 82294 70002 82350
rect 70058 82294 78970 82350
rect 79026 82294 79094 82350
rect 79150 82294 79218 82350
rect 79274 82294 79342 82350
rect 79398 82294 96970 82350
rect 97026 82294 97094 82350
rect 97150 82294 97218 82350
rect 97274 82294 97342 82350
rect 97398 82294 100598 82350
rect 100654 82294 100722 82350
rect 100778 82294 131318 82350
rect 131374 82294 131442 82350
rect 131498 82294 162038 82350
rect 162094 82294 162162 82350
rect 162218 82294 192758 82350
rect 192814 82294 192882 82350
rect 192938 82294 223478 82350
rect 223534 82294 223602 82350
rect 223658 82294 254198 82350
rect 254254 82294 254322 82350
rect 254378 82294 284918 82350
rect 284974 82294 285042 82350
rect 285098 82294 315638 82350
rect 315694 82294 315762 82350
rect 315818 82294 346358 82350
rect 346414 82294 346482 82350
rect 346538 82294 377078 82350
rect 377134 82294 377202 82350
rect 377258 82294 407798 82350
rect 407854 82294 407922 82350
rect 407978 82294 438518 82350
rect 438574 82294 438642 82350
rect 438698 82294 469238 82350
rect 469294 82294 469362 82350
rect 469418 82294 499958 82350
rect 500014 82294 500082 82350
rect 500138 82294 530678 82350
rect 530734 82294 530802 82350
rect 530858 82294 564970 82350
rect 565026 82294 565094 82350
rect 565150 82294 565218 82350
rect 565274 82294 565342 82350
rect 565398 82294 582970 82350
rect 583026 82294 583094 82350
rect 583150 82294 583218 82350
rect 583274 82294 583342 82350
rect 583398 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect -1916 82226 597980 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 6970 82226
rect 7026 82170 7094 82226
rect 7150 82170 7218 82226
rect 7274 82170 7342 82226
rect 7398 82170 24970 82226
rect 25026 82170 25094 82226
rect 25150 82170 25218 82226
rect 25274 82170 25342 82226
rect 25398 82170 42970 82226
rect 43026 82170 43094 82226
rect 43150 82170 43218 82226
rect 43274 82170 43342 82226
rect 43398 82170 60970 82226
rect 61026 82170 61094 82226
rect 61150 82170 61218 82226
rect 61274 82170 61342 82226
rect 61398 82170 69878 82226
rect 69934 82170 70002 82226
rect 70058 82170 78970 82226
rect 79026 82170 79094 82226
rect 79150 82170 79218 82226
rect 79274 82170 79342 82226
rect 79398 82170 96970 82226
rect 97026 82170 97094 82226
rect 97150 82170 97218 82226
rect 97274 82170 97342 82226
rect 97398 82170 100598 82226
rect 100654 82170 100722 82226
rect 100778 82170 131318 82226
rect 131374 82170 131442 82226
rect 131498 82170 162038 82226
rect 162094 82170 162162 82226
rect 162218 82170 192758 82226
rect 192814 82170 192882 82226
rect 192938 82170 223478 82226
rect 223534 82170 223602 82226
rect 223658 82170 254198 82226
rect 254254 82170 254322 82226
rect 254378 82170 284918 82226
rect 284974 82170 285042 82226
rect 285098 82170 315638 82226
rect 315694 82170 315762 82226
rect 315818 82170 346358 82226
rect 346414 82170 346482 82226
rect 346538 82170 377078 82226
rect 377134 82170 377202 82226
rect 377258 82170 407798 82226
rect 407854 82170 407922 82226
rect 407978 82170 438518 82226
rect 438574 82170 438642 82226
rect 438698 82170 469238 82226
rect 469294 82170 469362 82226
rect 469418 82170 499958 82226
rect 500014 82170 500082 82226
rect 500138 82170 530678 82226
rect 530734 82170 530802 82226
rect 530858 82170 564970 82226
rect 565026 82170 565094 82226
rect 565150 82170 565218 82226
rect 565274 82170 565342 82226
rect 565398 82170 582970 82226
rect 583026 82170 583094 82226
rect 583150 82170 583218 82226
rect 583274 82170 583342 82226
rect 583398 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect -1916 82102 597980 82170
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 6970 82102
rect 7026 82046 7094 82102
rect 7150 82046 7218 82102
rect 7274 82046 7342 82102
rect 7398 82046 24970 82102
rect 25026 82046 25094 82102
rect 25150 82046 25218 82102
rect 25274 82046 25342 82102
rect 25398 82046 42970 82102
rect 43026 82046 43094 82102
rect 43150 82046 43218 82102
rect 43274 82046 43342 82102
rect 43398 82046 60970 82102
rect 61026 82046 61094 82102
rect 61150 82046 61218 82102
rect 61274 82046 61342 82102
rect 61398 82046 69878 82102
rect 69934 82046 70002 82102
rect 70058 82046 78970 82102
rect 79026 82046 79094 82102
rect 79150 82046 79218 82102
rect 79274 82046 79342 82102
rect 79398 82046 96970 82102
rect 97026 82046 97094 82102
rect 97150 82046 97218 82102
rect 97274 82046 97342 82102
rect 97398 82046 100598 82102
rect 100654 82046 100722 82102
rect 100778 82046 131318 82102
rect 131374 82046 131442 82102
rect 131498 82046 162038 82102
rect 162094 82046 162162 82102
rect 162218 82046 192758 82102
rect 192814 82046 192882 82102
rect 192938 82046 223478 82102
rect 223534 82046 223602 82102
rect 223658 82046 254198 82102
rect 254254 82046 254322 82102
rect 254378 82046 284918 82102
rect 284974 82046 285042 82102
rect 285098 82046 315638 82102
rect 315694 82046 315762 82102
rect 315818 82046 346358 82102
rect 346414 82046 346482 82102
rect 346538 82046 377078 82102
rect 377134 82046 377202 82102
rect 377258 82046 407798 82102
rect 407854 82046 407922 82102
rect 407978 82046 438518 82102
rect 438574 82046 438642 82102
rect 438698 82046 469238 82102
rect 469294 82046 469362 82102
rect 469418 82046 499958 82102
rect 500014 82046 500082 82102
rect 500138 82046 530678 82102
rect 530734 82046 530802 82102
rect 530858 82046 564970 82102
rect 565026 82046 565094 82102
rect 565150 82046 565218 82102
rect 565274 82046 565342 82102
rect 565398 82046 582970 82102
rect 583026 82046 583094 82102
rect 583150 82046 583218 82102
rect 583274 82046 583342 82102
rect 583398 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect -1916 81978 597980 82046
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 6970 81978
rect 7026 81922 7094 81978
rect 7150 81922 7218 81978
rect 7274 81922 7342 81978
rect 7398 81922 24970 81978
rect 25026 81922 25094 81978
rect 25150 81922 25218 81978
rect 25274 81922 25342 81978
rect 25398 81922 42970 81978
rect 43026 81922 43094 81978
rect 43150 81922 43218 81978
rect 43274 81922 43342 81978
rect 43398 81922 60970 81978
rect 61026 81922 61094 81978
rect 61150 81922 61218 81978
rect 61274 81922 61342 81978
rect 61398 81922 69878 81978
rect 69934 81922 70002 81978
rect 70058 81922 78970 81978
rect 79026 81922 79094 81978
rect 79150 81922 79218 81978
rect 79274 81922 79342 81978
rect 79398 81922 96970 81978
rect 97026 81922 97094 81978
rect 97150 81922 97218 81978
rect 97274 81922 97342 81978
rect 97398 81922 100598 81978
rect 100654 81922 100722 81978
rect 100778 81922 131318 81978
rect 131374 81922 131442 81978
rect 131498 81922 162038 81978
rect 162094 81922 162162 81978
rect 162218 81922 192758 81978
rect 192814 81922 192882 81978
rect 192938 81922 223478 81978
rect 223534 81922 223602 81978
rect 223658 81922 254198 81978
rect 254254 81922 254322 81978
rect 254378 81922 284918 81978
rect 284974 81922 285042 81978
rect 285098 81922 315638 81978
rect 315694 81922 315762 81978
rect 315818 81922 346358 81978
rect 346414 81922 346482 81978
rect 346538 81922 377078 81978
rect 377134 81922 377202 81978
rect 377258 81922 407798 81978
rect 407854 81922 407922 81978
rect 407978 81922 438518 81978
rect 438574 81922 438642 81978
rect 438698 81922 469238 81978
rect 469294 81922 469362 81978
rect 469418 81922 499958 81978
rect 500014 81922 500082 81978
rect 500138 81922 530678 81978
rect 530734 81922 530802 81978
rect 530858 81922 564970 81978
rect 565026 81922 565094 81978
rect 565150 81922 565218 81978
rect 565274 81922 565342 81978
rect 565398 81922 582970 81978
rect 583026 81922 583094 81978
rect 583150 81922 583218 81978
rect 583274 81922 583342 81978
rect 583398 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect -1916 81826 597980 81922
rect -1916 76350 597980 76446
rect -1916 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 3250 76350
rect 3306 76294 3374 76350
rect 3430 76294 3498 76350
rect 3554 76294 3622 76350
rect 3678 76294 21250 76350
rect 21306 76294 21374 76350
rect 21430 76294 21498 76350
rect 21554 76294 21622 76350
rect 21678 76294 39250 76350
rect 39306 76294 39374 76350
rect 39430 76294 39498 76350
rect 39554 76294 39622 76350
rect 39678 76294 54518 76350
rect 54574 76294 54642 76350
rect 54698 76294 57250 76350
rect 57306 76294 57374 76350
rect 57430 76294 57498 76350
rect 57554 76294 57622 76350
rect 57678 76294 75250 76350
rect 75306 76294 75374 76350
rect 75430 76294 75498 76350
rect 75554 76294 75622 76350
rect 75678 76294 85238 76350
rect 85294 76294 85362 76350
rect 85418 76294 93250 76350
rect 93306 76294 93374 76350
rect 93430 76294 93498 76350
rect 93554 76294 93622 76350
rect 93678 76294 111250 76350
rect 111306 76294 111374 76350
rect 111430 76294 111498 76350
rect 111554 76294 111622 76350
rect 111678 76294 115958 76350
rect 116014 76294 116082 76350
rect 116138 76294 146678 76350
rect 146734 76294 146802 76350
rect 146858 76294 177398 76350
rect 177454 76294 177522 76350
rect 177578 76294 208118 76350
rect 208174 76294 208242 76350
rect 208298 76294 238838 76350
rect 238894 76294 238962 76350
rect 239018 76294 269558 76350
rect 269614 76294 269682 76350
rect 269738 76294 300278 76350
rect 300334 76294 300402 76350
rect 300458 76294 330998 76350
rect 331054 76294 331122 76350
rect 331178 76294 361718 76350
rect 361774 76294 361842 76350
rect 361898 76294 392438 76350
rect 392494 76294 392562 76350
rect 392618 76294 423158 76350
rect 423214 76294 423282 76350
rect 423338 76294 453878 76350
rect 453934 76294 454002 76350
rect 454058 76294 484598 76350
rect 484654 76294 484722 76350
rect 484778 76294 515318 76350
rect 515374 76294 515442 76350
rect 515498 76294 546038 76350
rect 546094 76294 546162 76350
rect 546218 76294 561250 76350
rect 561306 76294 561374 76350
rect 561430 76294 561498 76350
rect 561554 76294 561622 76350
rect 561678 76294 579250 76350
rect 579306 76294 579374 76350
rect 579430 76294 579498 76350
rect 579554 76294 579622 76350
rect 579678 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597980 76350
rect -1916 76226 597980 76294
rect -1916 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 3250 76226
rect 3306 76170 3374 76226
rect 3430 76170 3498 76226
rect 3554 76170 3622 76226
rect 3678 76170 21250 76226
rect 21306 76170 21374 76226
rect 21430 76170 21498 76226
rect 21554 76170 21622 76226
rect 21678 76170 39250 76226
rect 39306 76170 39374 76226
rect 39430 76170 39498 76226
rect 39554 76170 39622 76226
rect 39678 76170 54518 76226
rect 54574 76170 54642 76226
rect 54698 76170 57250 76226
rect 57306 76170 57374 76226
rect 57430 76170 57498 76226
rect 57554 76170 57622 76226
rect 57678 76170 75250 76226
rect 75306 76170 75374 76226
rect 75430 76170 75498 76226
rect 75554 76170 75622 76226
rect 75678 76170 85238 76226
rect 85294 76170 85362 76226
rect 85418 76170 93250 76226
rect 93306 76170 93374 76226
rect 93430 76170 93498 76226
rect 93554 76170 93622 76226
rect 93678 76170 111250 76226
rect 111306 76170 111374 76226
rect 111430 76170 111498 76226
rect 111554 76170 111622 76226
rect 111678 76170 115958 76226
rect 116014 76170 116082 76226
rect 116138 76170 146678 76226
rect 146734 76170 146802 76226
rect 146858 76170 177398 76226
rect 177454 76170 177522 76226
rect 177578 76170 208118 76226
rect 208174 76170 208242 76226
rect 208298 76170 238838 76226
rect 238894 76170 238962 76226
rect 239018 76170 269558 76226
rect 269614 76170 269682 76226
rect 269738 76170 300278 76226
rect 300334 76170 300402 76226
rect 300458 76170 330998 76226
rect 331054 76170 331122 76226
rect 331178 76170 361718 76226
rect 361774 76170 361842 76226
rect 361898 76170 392438 76226
rect 392494 76170 392562 76226
rect 392618 76170 423158 76226
rect 423214 76170 423282 76226
rect 423338 76170 453878 76226
rect 453934 76170 454002 76226
rect 454058 76170 484598 76226
rect 484654 76170 484722 76226
rect 484778 76170 515318 76226
rect 515374 76170 515442 76226
rect 515498 76170 546038 76226
rect 546094 76170 546162 76226
rect 546218 76170 561250 76226
rect 561306 76170 561374 76226
rect 561430 76170 561498 76226
rect 561554 76170 561622 76226
rect 561678 76170 579250 76226
rect 579306 76170 579374 76226
rect 579430 76170 579498 76226
rect 579554 76170 579622 76226
rect 579678 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597980 76226
rect -1916 76102 597980 76170
rect -1916 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 3250 76102
rect 3306 76046 3374 76102
rect 3430 76046 3498 76102
rect 3554 76046 3622 76102
rect 3678 76046 21250 76102
rect 21306 76046 21374 76102
rect 21430 76046 21498 76102
rect 21554 76046 21622 76102
rect 21678 76046 39250 76102
rect 39306 76046 39374 76102
rect 39430 76046 39498 76102
rect 39554 76046 39622 76102
rect 39678 76046 54518 76102
rect 54574 76046 54642 76102
rect 54698 76046 57250 76102
rect 57306 76046 57374 76102
rect 57430 76046 57498 76102
rect 57554 76046 57622 76102
rect 57678 76046 75250 76102
rect 75306 76046 75374 76102
rect 75430 76046 75498 76102
rect 75554 76046 75622 76102
rect 75678 76046 85238 76102
rect 85294 76046 85362 76102
rect 85418 76046 93250 76102
rect 93306 76046 93374 76102
rect 93430 76046 93498 76102
rect 93554 76046 93622 76102
rect 93678 76046 111250 76102
rect 111306 76046 111374 76102
rect 111430 76046 111498 76102
rect 111554 76046 111622 76102
rect 111678 76046 115958 76102
rect 116014 76046 116082 76102
rect 116138 76046 146678 76102
rect 146734 76046 146802 76102
rect 146858 76046 177398 76102
rect 177454 76046 177522 76102
rect 177578 76046 208118 76102
rect 208174 76046 208242 76102
rect 208298 76046 238838 76102
rect 238894 76046 238962 76102
rect 239018 76046 269558 76102
rect 269614 76046 269682 76102
rect 269738 76046 300278 76102
rect 300334 76046 300402 76102
rect 300458 76046 330998 76102
rect 331054 76046 331122 76102
rect 331178 76046 361718 76102
rect 361774 76046 361842 76102
rect 361898 76046 392438 76102
rect 392494 76046 392562 76102
rect 392618 76046 423158 76102
rect 423214 76046 423282 76102
rect 423338 76046 453878 76102
rect 453934 76046 454002 76102
rect 454058 76046 484598 76102
rect 484654 76046 484722 76102
rect 484778 76046 515318 76102
rect 515374 76046 515442 76102
rect 515498 76046 546038 76102
rect 546094 76046 546162 76102
rect 546218 76046 561250 76102
rect 561306 76046 561374 76102
rect 561430 76046 561498 76102
rect 561554 76046 561622 76102
rect 561678 76046 579250 76102
rect 579306 76046 579374 76102
rect 579430 76046 579498 76102
rect 579554 76046 579622 76102
rect 579678 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597980 76102
rect -1916 75978 597980 76046
rect -1916 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 3250 75978
rect 3306 75922 3374 75978
rect 3430 75922 3498 75978
rect 3554 75922 3622 75978
rect 3678 75922 21250 75978
rect 21306 75922 21374 75978
rect 21430 75922 21498 75978
rect 21554 75922 21622 75978
rect 21678 75922 39250 75978
rect 39306 75922 39374 75978
rect 39430 75922 39498 75978
rect 39554 75922 39622 75978
rect 39678 75922 54518 75978
rect 54574 75922 54642 75978
rect 54698 75922 57250 75978
rect 57306 75922 57374 75978
rect 57430 75922 57498 75978
rect 57554 75922 57622 75978
rect 57678 75922 75250 75978
rect 75306 75922 75374 75978
rect 75430 75922 75498 75978
rect 75554 75922 75622 75978
rect 75678 75922 85238 75978
rect 85294 75922 85362 75978
rect 85418 75922 93250 75978
rect 93306 75922 93374 75978
rect 93430 75922 93498 75978
rect 93554 75922 93622 75978
rect 93678 75922 111250 75978
rect 111306 75922 111374 75978
rect 111430 75922 111498 75978
rect 111554 75922 111622 75978
rect 111678 75922 115958 75978
rect 116014 75922 116082 75978
rect 116138 75922 146678 75978
rect 146734 75922 146802 75978
rect 146858 75922 177398 75978
rect 177454 75922 177522 75978
rect 177578 75922 208118 75978
rect 208174 75922 208242 75978
rect 208298 75922 238838 75978
rect 238894 75922 238962 75978
rect 239018 75922 269558 75978
rect 269614 75922 269682 75978
rect 269738 75922 300278 75978
rect 300334 75922 300402 75978
rect 300458 75922 330998 75978
rect 331054 75922 331122 75978
rect 331178 75922 361718 75978
rect 361774 75922 361842 75978
rect 361898 75922 392438 75978
rect 392494 75922 392562 75978
rect 392618 75922 423158 75978
rect 423214 75922 423282 75978
rect 423338 75922 453878 75978
rect 453934 75922 454002 75978
rect 454058 75922 484598 75978
rect 484654 75922 484722 75978
rect 484778 75922 515318 75978
rect 515374 75922 515442 75978
rect 515498 75922 546038 75978
rect 546094 75922 546162 75978
rect 546218 75922 561250 75978
rect 561306 75922 561374 75978
rect 561430 75922 561498 75978
rect 561554 75922 561622 75978
rect 561678 75922 579250 75978
rect 579306 75922 579374 75978
rect 579430 75922 579498 75978
rect 579554 75922 579622 75978
rect 579678 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597980 75978
rect -1916 75826 597980 75922
rect -1916 64350 597980 64446
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 6970 64350
rect 7026 64294 7094 64350
rect 7150 64294 7218 64350
rect 7274 64294 7342 64350
rect 7398 64294 24970 64350
rect 25026 64294 25094 64350
rect 25150 64294 25218 64350
rect 25274 64294 25342 64350
rect 25398 64294 42970 64350
rect 43026 64294 43094 64350
rect 43150 64294 43218 64350
rect 43274 64294 43342 64350
rect 43398 64294 60970 64350
rect 61026 64294 61094 64350
rect 61150 64294 61218 64350
rect 61274 64294 61342 64350
rect 61398 64294 69878 64350
rect 69934 64294 70002 64350
rect 70058 64294 78970 64350
rect 79026 64294 79094 64350
rect 79150 64294 79218 64350
rect 79274 64294 79342 64350
rect 79398 64294 96970 64350
rect 97026 64294 97094 64350
rect 97150 64294 97218 64350
rect 97274 64294 97342 64350
rect 97398 64294 100598 64350
rect 100654 64294 100722 64350
rect 100778 64294 131318 64350
rect 131374 64294 131442 64350
rect 131498 64294 162038 64350
rect 162094 64294 162162 64350
rect 162218 64294 192758 64350
rect 192814 64294 192882 64350
rect 192938 64294 223478 64350
rect 223534 64294 223602 64350
rect 223658 64294 254198 64350
rect 254254 64294 254322 64350
rect 254378 64294 284918 64350
rect 284974 64294 285042 64350
rect 285098 64294 315638 64350
rect 315694 64294 315762 64350
rect 315818 64294 346358 64350
rect 346414 64294 346482 64350
rect 346538 64294 377078 64350
rect 377134 64294 377202 64350
rect 377258 64294 407798 64350
rect 407854 64294 407922 64350
rect 407978 64294 438518 64350
rect 438574 64294 438642 64350
rect 438698 64294 469238 64350
rect 469294 64294 469362 64350
rect 469418 64294 499958 64350
rect 500014 64294 500082 64350
rect 500138 64294 530678 64350
rect 530734 64294 530802 64350
rect 530858 64294 564970 64350
rect 565026 64294 565094 64350
rect 565150 64294 565218 64350
rect 565274 64294 565342 64350
rect 565398 64294 582970 64350
rect 583026 64294 583094 64350
rect 583150 64294 583218 64350
rect 583274 64294 583342 64350
rect 583398 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect -1916 64226 597980 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 6970 64226
rect 7026 64170 7094 64226
rect 7150 64170 7218 64226
rect 7274 64170 7342 64226
rect 7398 64170 24970 64226
rect 25026 64170 25094 64226
rect 25150 64170 25218 64226
rect 25274 64170 25342 64226
rect 25398 64170 42970 64226
rect 43026 64170 43094 64226
rect 43150 64170 43218 64226
rect 43274 64170 43342 64226
rect 43398 64170 60970 64226
rect 61026 64170 61094 64226
rect 61150 64170 61218 64226
rect 61274 64170 61342 64226
rect 61398 64170 69878 64226
rect 69934 64170 70002 64226
rect 70058 64170 78970 64226
rect 79026 64170 79094 64226
rect 79150 64170 79218 64226
rect 79274 64170 79342 64226
rect 79398 64170 96970 64226
rect 97026 64170 97094 64226
rect 97150 64170 97218 64226
rect 97274 64170 97342 64226
rect 97398 64170 100598 64226
rect 100654 64170 100722 64226
rect 100778 64170 131318 64226
rect 131374 64170 131442 64226
rect 131498 64170 162038 64226
rect 162094 64170 162162 64226
rect 162218 64170 192758 64226
rect 192814 64170 192882 64226
rect 192938 64170 223478 64226
rect 223534 64170 223602 64226
rect 223658 64170 254198 64226
rect 254254 64170 254322 64226
rect 254378 64170 284918 64226
rect 284974 64170 285042 64226
rect 285098 64170 315638 64226
rect 315694 64170 315762 64226
rect 315818 64170 346358 64226
rect 346414 64170 346482 64226
rect 346538 64170 377078 64226
rect 377134 64170 377202 64226
rect 377258 64170 407798 64226
rect 407854 64170 407922 64226
rect 407978 64170 438518 64226
rect 438574 64170 438642 64226
rect 438698 64170 469238 64226
rect 469294 64170 469362 64226
rect 469418 64170 499958 64226
rect 500014 64170 500082 64226
rect 500138 64170 530678 64226
rect 530734 64170 530802 64226
rect 530858 64170 564970 64226
rect 565026 64170 565094 64226
rect 565150 64170 565218 64226
rect 565274 64170 565342 64226
rect 565398 64170 582970 64226
rect 583026 64170 583094 64226
rect 583150 64170 583218 64226
rect 583274 64170 583342 64226
rect 583398 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect -1916 64102 597980 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 6970 64102
rect 7026 64046 7094 64102
rect 7150 64046 7218 64102
rect 7274 64046 7342 64102
rect 7398 64046 24970 64102
rect 25026 64046 25094 64102
rect 25150 64046 25218 64102
rect 25274 64046 25342 64102
rect 25398 64046 42970 64102
rect 43026 64046 43094 64102
rect 43150 64046 43218 64102
rect 43274 64046 43342 64102
rect 43398 64046 60970 64102
rect 61026 64046 61094 64102
rect 61150 64046 61218 64102
rect 61274 64046 61342 64102
rect 61398 64046 69878 64102
rect 69934 64046 70002 64102
rect 70058 64046 78970 64102
rect 79026 64046 79094 64102
rect 79150 64046 79218 64102
rect 79274 64046 79342 64102
rect 79398 64046 96970 64102
rect 97026 64046 97094 64102
rect 97150 64046 97218 64102
rect 97274 64046 97342 64102
rect 97398 64046 100598 64102
rect 100654 64046 100722 64102
rect 100778 64046 131318 64102
rect 131374 64046 131442 64102
rect 131498 64046 162038 64102
rect 162094 64046 162162 64102
rect 162218 64046 192758 64102
rect 192814 64046 192882 64102
rect 192938 64046 223478 64102
rect 223534 64046 223602 64102
rect 223658 64046 254198 64102
rect 254254 64046 254322 64102
rect 254378 64046 284918 64102
rect 284974 64046 285042 64102
rect 285098 64046 315638 64102
rect 315694 64046 315762 64102
rect 315818 64046 346358 64102
rect 346414 64046 346482 64102
rect 346538 64046 377078 64102
rect 377134 64046 377202 64102
rect 377258 64046 407798 64102
rect 407854 64046 407922 64102
rect 407978 64046 438518 64102
rect 438574 64046 438642 64102
rect 438698 64046 469238 64102
rect 469294 64046 469362 64102
rect 469418 64046 499958 64102
rect 500014 64046 500082 64102
rect 500138 64046 530678 64102
rect 530734 64046 530802 64102
rect 530858 64046 564970 64102
rect 565026 64046 565094 64102
rect 565150 64046 565218 64102
rect 565274 64046 565342 64102
rect 565398 64046 582970 64102
rect 583026 64046 583094 64102
rect 583150 64046 583218 64102
rect 583274 64046 583342 64102
rect 583398 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect -1916 63978 597980 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 6970 63978
rect 7026 63922 7094 63978
rect 7150 63922 7218 63978
rect 7274 63922 7342 63978
rect 7398 63922 24970 63978
rect 25026 63922 25094 63978
rect 25150 63922 25218 63978
rect 25274 63922 25342 63978
rect 25398 63922 42970 63978
rect 43026 63922 43094 63978
rect 43150 63922 43218 63978
rect 43274 63922 43342 63978
rect 43398 63922 60970 63978
rect 61026 63922 61094 63978
rect 61150 63922 61218 63978
rect 61274 63922 61342 63978
rect 61398 63922 69878 63978
rect 69934 63922 70002 63978
rect 70058 63922 78970 63978
rect 79026 63922 79094 63978
rect 79150 63922 79218 63978
rect 79274 63922 79342 63978
rect 79398 63922 96970 63978
rect 97026 63922 97094 63978
rect 97150 63922 97218 63978
rect 97274 63922 97342 63978
rect 97398 63922 100598 63978
rect 100654 63922 100722 63978
rect 100778 63922 131318 63978
rect 131374 63922 131442 63978
rect 131498 63922 162038 63978
rect 162094 63922 162162 63978
rect 162218 63922 192758 63978
rect 192814 63922 192882 63978
rect 192938 63922 223478 63978
rect 223534 63922 223602 63978
rect 223658 63922 254198 63978
rect 254254 63922 254322 63978
rect 254378 63922 284918 63978
rect 284974 63922 285042 63978
rect 285098 63922 315638 63978
rect 315694 63922 315762 63978
rect 315818 63922 346358 63978
rect 346414 63922 346482 63978
rect 346538 63922 377078 63978
rect 377134 63922 377202 63978
rect 377258 63922 407798 63978
rect 407854 63922 407922 63978
rect 407978 63922 438518 63978
rect 438574 63922 438642 63978
rect 438698 63922 469238 63978
rect 469294 63922 469362 63978
rect 469418 63922 499958 63978
rect 500014 63922 500082 63978
rect 500138 63922 530678 63978
rect 530734 63922 530802 63978
rect 530858 63922 564970 63978
rect 565026 63922 565094 63978
rect 565150 63922 565218 63978
rect 565274 63922 565342 63978
rect 565398 63922 582970 63978
rect 583026 63922 583094 63978
rect 583150 63922 583218 63978
rect 583274 63922 583342 63978
rect 583398 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect -1916 63826 597980 63922
rect -1916 58350 597980 58446
rect -1916 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 3250 58350
rect 3306 58294 3374 58350
rect 3430 58294 3498 58350
rect 3554 58294 3622 58350
rect 3678 58294 21250 58350
rect 21306 58294 21374 58350
rect 21430 58294 21498 58350
rect 21554 58294 21622 58350
rect 21678 58294 39250 58350
rect 39306 58294 39374 58350
rect 39430 58294 39498 58350
rect 39554 58294 39622 58350
rect 39678 58294 54518 58350
rect 54574 58294 54642 58350
rect 54698 58294 57250 58350
rect 57306 58294 57374 58350
rect 57430 58294 57498 58350
rect 57554 58294 57622 58350
rect 57678 58294 75250 58350
rect 75306 58294 75374 58350
rect 75430 58294 75498 58350
rect 75554 58294 75622 58350
rect 75678 58294 85238 58350
rect 85294 58294 85362 58350
rect 85418 58294 93250 58350
rect 93306 58294 93374 58350
rect 93430 58294 93498 58350
rect 93554 58294 93622 58350
rect 93678 58294 111250 58350
rect 111306 58294 111374 58350
rect 111430 58294 111498 58350
rect 111554 58294 111622 58350
rect 111678 58294 115958 58350
rect 116014 58294 116082 58350
rect 116138 58294 146678 58350
rect 146734 58294 146802 58350
rect 146858 58294 177398 58350
rect 177454 58294 177522 58350
rect 177578 58294 208118 58350
rect 208174 58294 208242 58350
rect 208298 58294 238838 58350
rect 238894 58294 238962 58350
rect 239018 58294 269558 58350
rect 269614 58294 269682 58350
rect 269738 58294 300278 58350
rect 300334 58294 300402 58350
rect 300458 58294 330998 58350
rect 331054 58294 331122 58350
rect 331178 58294 361718 58350
rect 361774 58294 361842 58350
rect 361898 58294 392438 58350
rect 392494 58294 392562 58350
rect 392618 58294 423158 58350
rect 423214 58294 423282 58350
rect 423338 58294 453878 58350
rect 453934 58294 454002 58350
rect 454058 58294 484598 58350
rect 484654 58294 484722 58350
rect 484778 58294 515318 58350
rect 515374 58294 515442 58350
rect 515498 58294 546038 58350
rect 546094 58294 546162 58350
rect 546218 58294 561250 58350
rect 561306 58294 561374 58350
rect 561430 58294 561498 58350
rect 561554 58294 561622 58350
rect 561678 58294 579250 58350
rect 579306 58294 579374 58350
rect 579430 58294 579498 58350
rect 579554 58294 579622 58350
rect 579678 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597980 58350
rect -1916 58226 597980 58294
rect -1916 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 3250 58226
rect 3306 58170 3374 58226
rect 3430 58170 3498 58226
rect 3554 58170 3622 58226
rect 3678 58170 21250 58226
rect 21306 58170 21374 58226
rect 21430 58170 21498 58226
rect 21554 58170 21622 58226
rect 21678 58170 39250 58226
rect 39306 58170 39374 58226
rect 39430 58170 39498 58226
rect 39554 58170 39622 58226
rect 39678 58170 54518 58226
rect 54574 58170 54642 58226
rect 54698 58170 57250 58226
rect 57306 58170 57374 58226
rect 57430 58170 57498 58226
rect 57554 58170 57622 58226
rect 57678 58170 75250 58226
rect 75306 58170 75374 58226
rect 75430 58170 75498 58226
rect 75554 58170 75622 58226
rect 75678 58170 85238 58226
rect 85294 58170 85362 58226
rect 85418 58170 93250 58226
rect 93306 58170 93374 58226
rect 93430 58170 93498 58226
rect 93554 58170 93622 58226
rect 93678 58170 111250 58226
rect 111306 58170 111374 58226
rect 111430 58170 111498 58226
rect 111554 58170 111622 58226
rect 111678 58170 115958 58226
rect 116014 58170 116082 58226
rect 116138 58170 146678 58226
rect 146734 58170 146802 58226
rect 146858 58170 177398 58226
rect 177454 58170 177522 58226
rect 177578 58170 208118 58226
rect 208174 58170 208242 58226
rect 208298 58170 238838 58226
rect 238894 58170 238962 58226
rect 239018 58170 269558 58226
rect 269614 58170 269682 58226
rect 269738 58170 300278 58226
rect 300334 58170 300402 58226
rect 300458 58170 330998 58226
rect 331054 58170 331122 58226
rect 331178 58170 361718 58226
rect 361774 58170 361842 58226
rect 361898 58170 392438 58226
rect 392494 58170 392562 58226
rect 392618 58170 423158 58226
rect 423214 58170 423282 58226
rect 423338 58170 453878 58226
rect 453934 58170 454002 58226
rect 454058 58170 484598 58226
rect 484654 58170 484722 58226
rect 484778 58170 515318 58226
rect 515374 58170 515442 58226
rect 515498 58170 546038 58226
rect 546094 58170 546162 58226
rect 546218 58170 561250 58226
rect 561306 58170 561374 58226
rect 561430 58170 561498 58226
rect 561554 58170 561622 58226
rect 561678 58170 579250 58226
rect 579306 58170 579374 58226
rect 579430 58170 579498 58226
rect 579554 58170 579622 58226
rect 579678 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597980 58226
rect -1916 58102 597980 58170
rect -1916 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 3250 58102
rect 3306 58046 3374 58102
rect 3430 58046 3498 58102
rect 3554 58046 3622 58102
rect 3678 58046 21250 58102
rect 21306 58046 21374 58102
rect 21430 58046 21498 58102
rect 21554 58046 21622 58102
rect 21678 58046 39250 58102
rect 39306 58046 39374 58102
rect 39430 58046 39498 58102
rect 39554 58046 39622 58102
rect 39678 58046 54518 58102
rect 54574 58046 54642 58102
rect 54698 58046 57250 58102
rect 57306 58046 57374 58102
rect 57430 58046 57498 58102
rect 57554 58046 57622 58102
rect 57678 58046 75250 58102
rect 75306 58046 75374 58102
rect 75430 58046 75498 58102
rect 75554 58046 75622 58102
rect 75678 58046 85238 58102
rect 85294 58046 85362 58102
rect 85418 58046 93250 58102
rect 93306 58046 93374 58102
rect 93430 58046 93498 58102
rect 93554 58046 93622 58102
rect 93678 58046 111250 58102
rect 111306 58046 111374 58102
rect 111430 58046 111498 58102
rect 111554 58046 111622 58102
rect 111678 58046 115958 58102
rect 116014 58046 116082 58102
rect 116138 58046 146678 58102
rect 146734 58046 146802 58102
rect 146858 58046 177398 58102
rect 177454 58046 177522 58102
rect 177578 58046 208118 58102
rect 208174 58046 208242 58102
rect 208298 58046 238838 58102
rect 238894 58046 238962 58102
rect 239018 58046 269558 58102
rect 269614 58046 269682 58102
rect 269738 58046 300278 58102
rect 300334 58046 300402 58102
rect 300458 58046 330998 58102
rect 331054 58046 331122 58102
rect 331178 58046 361718 58102
rect 361774 58046 361842 58102
rect 361898 58046 392438 58102
rect 392494 58046 392562 58102
rect 392618 58046 423158 58102
rect 423214 58046 423282 58102
rect 423338 58046 453878 58102
rect 453934 58046 454002 58102
rect 454058 58046 484598 58102
rect 484654 58046 484722 58102
rect 484778 58046 515318 58102
rect 515374 58046 515442 58102
rect 515498 58046 546038 58102
rect 546094 58046 546162 58102
rect 546218 58046 561250 58102
rect 561306 58046 561374 58102
rect 561430 58046 561498 58102
rect 561554 58046 561622 58102
rect 561678 58046 579250 58102
rect 579306 58046 579374 58102
rect 579430 58046 579498 58102
rect 579554 58046 579622 58102
rect 579678 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597980 58102
rect -1916 57978 597980 58046
rect -1916 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 3250 57978
rect 3306 57922 3374 57978
rect 3430 57922 3498 57978
rect 3554 57922 3622 57978
rect 3678 57922 21250 57978
rect 21306 57922 21374 57978
rect 21430 57922 21498 57978
rect 21554 57922 21622 57978
rect 21678 57922 39250 57978
rect 39306 57922 39374 57978
rect 39430 57922 39498 57978
rect 39554 57922 39622 57978
rect 39678 57922 54518 57978
rect 54574 57922 54642 57978
rect 54698 57922 57250 57978
rect 57306 57922 57374 57978
rect 57430 57922 57498 57978
rect 57554 57922 57622 57978
rect 57678 57922 75250 57978
rect 75306 57922 75374 57978
rect 75430 57922 75498 57978
rect 75554 57922 75622 57978
rect 75678 57922 85238 57978
rect 85294 57922 85362 57978
rect 85418 57922 93250 57978
rect 93306 57922 93374 57978
rect 93430 57922 93498 57978
rect 93554 57922 93622 57978
rect 93678 57922 111250 57978
rect 111306 57922 111374 57978
rect 111430 57922 111498 57978
rect 111554 57922 111622 57978
rect 111678 57922 115958 57978
rect 116014 57922 116082 57978
rect 116138 57922 146678 57978
rect 146734 57922 146802 57978
rect 146858 57922 177398 57978
rect 177454 57922 177522 57978
rect 177578 57922 208118 57978
rect 208174 57922 208242 57978
rect 208298 57922 238838 57978
rect 238894 57922 238962 57978
rect 239018 57922 269558 57978
rect 269614 57922 269682 57978
rect 269738 57922 300278 57978
rect 300334 57922 300402 57978
rect 300458 57922 330998 57978
rect 331054 57922 331122 57978
rect 331178 57922 361718 57978
rect 361774 57922 361842 57978
rect 361898 57922 392438 57978
rect 392494 57922 392562 57978
rect 392618 57922 423158 57978
rect 423214 57922 423282 57978
rect 423338 57922 453878 57978
rect 453934 57922 454002 57978
rect 454058 57922 484598 57978
rect 484654 57922 484722 57978
rect 484778 57922 515318 57978
rect 515374 57922 515442 57978
rect 515498 57922 546038 57978
rect 546094 57922 546162 57978
rect 546218 57922 561250 57978
rect 561306 57922 561374 57978
rect 561430 57922 561498 57978
rect 561554 57922 561622 57978
rect 561678 57922 579250 57978
rect 579306 57922 579374 57978
rect 579430 57922 579498 57978
rect 579554 57922 579622 57978
rect 579678 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597980 57978
rect -1916 57826 597980 57922
rect -1916 46350 597980 46446
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 6970 46350
rect 7026 46294 7094 46350
rect 7150 46294 7218 46350
rect 7274 46294 7342 46350
rect 7398 46294 24970 46350
rect 25026 46294 25094 46350
rect 25150 46294 25218 46350
rect 25274 46294 25342 46350
rect 25398 46294 42970 46350
rect 43026 46294 43094 46350
rect 43150 46294 43218 46350
rect 43274 46294 43342 46350
rect 43398 46294 60970 46350
rect 61026 46294 61094 46350
rect 61150 46294 61218 46350
rect 61274 46294 61342 46350
rect 61398 46294 69878 46350
rect 69934 46294 70002 46350
rect 70058 46294 78970 46350
rect 79026 46294 79094 46350
rect 79150 46294 79218 46350
rect 79274 46294 79342 46350
rect 79398 46294 96970 46350
rect 97026 46294 97094 46350
rect 97150 46294 97218 46350
rect 97274 46294 97342 46350
rect 97398 46294 100598 46350
rect 100654 46294 100722 46350
rect 100778 46294 131318 46350
rect 131374 46294 131442 46350
rect 131498 46294 162038 46350
rect 162094 46294 162162 46350
rect 162218 46294 192758 46350
rect 192814 46294 192882 46350
rect 192938 46294 223478 46350
rect 223534 46294 223602 46350
rect 223658 46294 254198 46350
rect 254254 46294 254322 46350
rect 254378 46294 284918 46350
rect 284974 46294 285042 46350
rect 285098 46294 315638 46350
rect 315694 46294 315762 46350
rect 315818 46294 346358 46350
rect 346414 46294 346482 46350
rect 346538 46294 377078 46350
rect 377134 46294 377202 46350
rect 377258 46294 407798 46350
rect 407854 46294 407922 46350
rect 407978 46294 438518 46350
rect 438574 46294 438642 46350
rect 438698 46294 469238 46350
rect 469294 46294 469362 46350
rect 469418 46294 499958 46350
rect 500014 46294 500082 46350
rect 500138 46294 530678 46350
rect 530734 46294 530802 46350
rect 530858 46294 564970 46350
rect 565026 46294 565094 46350
rect 565150 46294 565218 46350
rect 565274 46294 565342 46350
rect 565398 46294 582970 46350
rect 583026 46294 583094 46350
rect 583150 46294 583218 46350
rect 583274 46294 583342 46350
rect 583398 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect -1916 46226 597980 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 6970 46226
rect 7026 46170 7094 46226
rect 7150 46170 7218 46226
rect 7274 46170 7342 46226
rect 7398 46170 24970 46226
rect 25026 46170 25094 46226
rect 25150 46170 25218 46226
rect 25274 46170 25342 46226
rect 25398 46170 42970 46226
rect 43026 46170 43094 46226
rect 43150 46170 43218 46226
rect 43274 46170 43342 46226
rect 43398 46170 60970 46226
rect 61026 46170 61094 46226
rect 61150 46170 61218 46226
rect 61274 46170 61342 46226
rect 61398 46170 69878 46226
rect 69934 46170 70002 46226
rect 70058 46170 78970 46226
rect 79026 46170 79094 46226
rect 79150 46170 79218 46226
rect 79274 46170 79342 46226
rect 79398 46170 96970 46226
rect 97026 46170 97094 46226
rect 97150 46170 97218 46226
rect 97274 46170 97342 46226
rect 97398 46170 100598 46226
rect 100654 46170 100722 46226
rect 100778 46170 131318 46226
rect 131374 46170 131442 46226
rect 131498 46170 162038 46226
rect 162094 46170 162162 46226
rect 162218 46170 192758 46226
rect 192814 46170 192882 46226
rect 192938 46170 223478 46226
rect 223534 46170 223602 46226
rect 223658 46170 254198 46226
rect 254254 46170 254322 46226
rect 254378 46170 284918 46226
rect 284974 46170 285042 46226
rect 285098 46170 315638 46226
rect 315694 46170 315762 46226
rect 315818 46170 346358 46226
rect 346414 46170 346482 46226
rect 346538 46170 377078 46226
rect 377134 46170 377202 46226
rect 377258 46170 407798 46226
rect 407854 46170 407922 46226
rect 407978 46170 438518 46226
rect 438574 46170 438642 46226
rect 438698 46170 469238 46226
rect 469294 46170 469362 46226
rect 469418 46170 499958 46226
rect 500014 46170 500082 46226
rect 500138 46170 530678 46226
rect 530734 46170 530802 46226
rect 530858 46170 564970 46226
rect 565026 46170 565094 46226
rect 565150 46170 565218 46226
rect 565274 46170 565342 46226
rect 565398 46170 582970 46226
rect 583026 46170 583094 46226
rect 583150 46170 583218 46226
rect 583274 46170 583342 46226
rect 583398 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect -1916 46102 597980 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 6970 46102
rect 7026 46046 7094 46102
rect 7150 46046 7218 46102
rect 7274 46046 7342 46102
rect 7398 46046 24970 46102
rect 25026 46046 25094 46102
rect 25150 46046 25218 46102
rect 25274 46046 25342 46102
rect 25398 46046 42970 46102
rect 43026 46046 43094 46102
rect 43150 46046 43218 46102
rect 43274 46046 43342 46102
rect 43398 46046 60970 46102
rect 61026 46046 61094 46102
rect 61150 46046 61218 46102
rect 61274 46046 61342 46102
rect 61398 46046 69878 46102
rect 69934 46046 70002 46102
rect 70058 46046 78970 46102
rect 79026 46046 79094 46102
rect 79150 46046 79218 46102
rect 79274 46046 79342 46102
rect 79398 46046 96970 46102
rect 97026 46046 97094 46102
rect 97150 46046 97218 46102
rect 97274 46046 97342 46102
rect 97398 46046 100598 46102
rect 100654 46046 100722 46102
rect 100778 46046 131318 46102
rect 131374 46046 131442 46102
rect 131498 46046 162038 46102
rect 162094 46046 162162 46102
rect 162218 46046 192758 46102
rect 192814 46046 192882 46102
rect 192938 46046 223478 46102
rect 223534 46046 223602 46102
rect 223658 46046 254198 46102
rect 254254 46046 254322 46102
rect 254378 46046 284918 46102
rect 284974 46046 285042 46102
rect 285098 46046 315638 46102
rect 315694 46046 315762 46102
rect 315818 46046 346358 46102
rect 346414 46046 346482 46102
rect 346538 46046 377078 46102
rect 377134 46046 377202 46102
rect 377258 46046 407798 46102
rect 407854 46046 407922 46102
rect 407978 46046 438518 46102
rect 438574 46046 438642 46102
rect 438698 46046 469238 46102
rect 469294 46046 469362 46102
rect 469418 46046 499958 46102
rect 500014 46046 500082 46102
rect 500138 46046 530678 46102
rect 530734 46046 530802 46102
rect 530858 46046 564970 46102
rect 565026 46046 565094 46102
rect 565150 46046 565218 46102
rect 565274 46046 565342 46102
rect 565398 46046 582970 46102
rect 583026 46046 583094 46102
rect 583150 46046 583218 46102
rect 583274 46046 583342 46102
rect 583398 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect -1916 45978 597980 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 6970 45978
rect 7026 45922 7094 45978
rect 7150 45922 7218 45978
rect 7274 45922 7342 45978
rect 7398 45922 24970 45978
rect 25026 45922 25094 45978
rect 25150 45922 25218 45978
rect 25274 45922 25342 45978
rect 25398 45922 42970 45978
rect 43026 45922 43094 45978
rect 43150 45922 43218 45978
rect 43274 45922 43342 45978
rect 43398 45922 60970 45978
rect 61026 45922 61094 45978
rect 61150 45922 61218 45978
rect 61274 45922 61342 45978
rect 61398 45922 69878 45978
rect 69934 45922 70002 45978
rect 70058 45922 78970 45978
rect 79026 45922 79094 45978
rect 79150 45922 79218 45978
rect 79274 45922 79342 45978
rect 79398 45922 96970 45978
rect 97026 45922 97094 45978
rect 97150 45922 97218 45978
rect 97274 45922 97342 45978
rect 97398 45922 100598 45978
rect 100654 45922 100722 45978
rect 100778 45922 131318 45978
rect 131374 45922 131442 45978
rect 131498 45922 162038 45978
rect 162094 45922 162162 45978
rect 162218 45922 192758 45978
rect 192814 45922 192882 45978
rect 192938 45922 223478 45978
rect 223534 45922 223602 45978
rect 223658 45922 254198 45978
rect 254254 45922 254322 45978
rect 254378 45922 284918 45978
rect 284974 45922 285042 45978
rect 285098 45922 315638 45978
rect 315694 45922 315762 45978
rect 315818 45922 346358 45978
rect 346414 45922 346482 45978
rect 346538 45922 377078 45978
rect 377134 45922 377202 45978
rect 377258 45922 407798 45978
rect 407854 45922 407922 45978
rect 407978 45922 438518 45978
rect 438574 45922 438642 45978
rect 438698 45922 469238 45978
rect 469294 45922 469362 45978
rect 469418 45922 499958 45978
rect 500014 45922 500082 45978
rect 500138 45922 530678 45978
rect 530734 45922 530802 45978
rect 530858 45922 564970 45978
rect 565026 45922 565094 45978
rect 565150 45922 565218 45978
rect 565274 45922 565342 45978
rect 565398 45922 582970 45978
rect 583026 45922 583094 45978
rect 583150 45922 583218 45978
rect 583274 45922 583342 45978
rect 583398 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect -1916 45826 597980 45922
rect -1916 40350 597980 40446
rect -1916 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 3250 40350
rect 3306 40294 3374 40350
rect 3430 40294 3498 40350
rect 3554 40294 3622 40350
rect 3678 40294 21250 40350
rect 21306 40294 21374 40350
rect 21430 40294 21498 40350
rect 21554 40294 21622 40350
rect 21678 40294 39250 40350
rect 39306 40294 39374 40350
rect 39430 40294 39498 40350
rect 39554 40294 39622 40350
rect 39678 40294 54518 40350
rect 54574 40294 54642 40350
rect 54698 40294 57250 40350
rect 57306 40294 57374 40350
rect 57430 40294 57498 40350
rect 57554 40294 57622 40350
rect 57678 40294 75250 40350
rect 75306 40294 75374 40350
rect 75430 40294 75498 40350
rect 75554 40294 75622 40350
rect 75678 40294 85238 40350
rect 85294 40294 85362 40350
rect 85418 40294 93250 40350
rect 93306 40294 93374 40350
rect 93430 40294 93498 40350
rect 93554 40294 93622 40350
rect 93678 40294 111250 40350
rect 111306 40294 111374 40350
rect 111430 40294 111498 40350
rect 111554 40294 111622 40350
rect 111678 40294 115958 40350
rect 116014 40294 116082 40350
rect 116138 40294 146678 40350
rect 146734 40294 146802 40350
rect 146858 40294 177398 40350
rect 177454 40294 177522 40350
rect 177578 40294 208118 40350
rect 208174 40294 208242 40350
rect 208298 40294 238838 40350
rect 238894 40294 238962 40350
rect 239018 40294 269558 40350
rect 269614 40294 269682 40350
rect 269738 40294 300278 40350
rect 300334 40294 300402 40350
rect 300458 40294 330998 40350
rect 331054 40294 331122 40350
rect 331178 40294 361718 40350
rect 361774 40294 361842 40350
rect 361898 40294 392438 40350
rect 392494 40294 392562 40350
rect 392618 40294 423158 40350
rect 423214 40294 423282 40350
rect 423338 40294 453878 40350
rect 453934 40294 454002 40350
rect 454058 40294 484598 40350
rect 484654 40294 484722 40350
rect 484778 40294 515318 40350
rect 515374 40294 515442 40350
rect 515498 40294 546038 40350
rect 546094 40294 546162 40350
rect 546218 40294 561250 40350
rect 561306 40294 561374 40350
rect 561430 40294 561498 40350
rect 561554 40294 561622 40350
rect 561678 40294 579250 40350
rect 579306 40294 579374 40350
rect 579430 40294 579498 40350
rect 579554 40294 579622 40350
rect 579678 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597980 40350
rect -1916 40226 597980 40294
rect -1916 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 3250 40226
rect 3306 40170 3374 40226
rect 3430 40170 3498 40226
rect 3554 40170 3622 40226
rect 3678 40170 21250 40226
rect 21306 40170 21374 40226
rect 21430 40170 21498 40226
rect 21554 40170 21622 40226
rect 21678 40170 39250 40226
rect 39306 40170 39374 40226
rect 39430 40170 39498 40226
rect 39554 40170 39622 40226
rect 39678 40170 54518 40226
rect 54574 40170 54642 40226
rect 54698 40170 57250 40226
rect 57306 40170 57374 40226
rect 57430 40170 57498 40226
rect 57554 40170 57622 40226
rect 57678 40170 75250 40226
rect 75306 40170 75374 40226
rect 75430 40170 75498 40226
rect 75554 40170 75622 40226
rect 75678 40170 85238 40226
rect 85294 40170 85362 40226
rect 85418 40170 93250 40226
rect 93306 40170 93374 40226
rect 93430 40170 93498 40226
rect 93554 40170 93622 40226
rect 93678 40170 111250 40226
rect 111306 40170 111374 40226
rect 111430 40170 111498 40226
rect 111554 40170 111622 40226
rect 111678 40170 115958 40226
rect 116014 40170 116082 40226
rect 116138 40170 146678 40226
rect 146734 40170 146802 40226
rect 146858 40170 177398 40226
rect 177454 40170 177522 40226
rect 177578 40170 208118 40226
rect 208174 40170 208242 40226
rect 208298 40170 238838 40226
rect 238894 40170 238962 40226
rect 239018 40170 269558 40226
rect 269614 40170 269682 40226
rect 269738 40170 300278 40226
rect 300334 40170 300402 40226
rect 300458 40170 330998 40226
rect 331054 40170 331122 40226
rect 331178 40170 361718 40226
rect 361774 40170 361842 40226
rect 361898 40170 392438 40226
rect 392494 40170 392562 40226
rect 392618 40170 423158 40226
rect 423214 40170 423282 40226
rect 423338 40170 453878 40226
rect 453934 40170 454002 40226
rect 454058 40170 484598 40226
rect 484654 40170 484722 40226
rect 484778 40170 515318 40226
rect 515374 40170 515442 40226
rect 515498 40170 546038 40226
rect 546094 40170 546162 40226
rect 546218 40170 561250 40226
rect 561306 40170 561374 40226
rect 561430 40170 561498 40226
rect 561554 40170 561622 40226
rect 561678 40170 579250 40226
rect 579306 40170 579374 40226
rect 579430 40170 579498 40226
rect 579554 40170 579622 40226
rect 579678 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597980 40226
rect -1916 40102 597980 40170
rect -1916 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 3250 40102
rect 3306 40046 3374 40102
rect 3430 40046 3498 40102
rect 3554 40046 3622 40102
rect 3678 40046 21250 40102
rect 21306 40046 21374 40102
rect 21430 40046 21498 40102
rect 21554 40046 21622 40102
rect 21678 40046 39250 40102
rect 39306 40046 39374 40102
rect 39430 40046 39498 40102
rect 39554 40046 39622 40102
rect 39678 40046 54518 40102
rect 54574 40046 54642 40102
rect 54698 40046 57250 40102
rect 57306 40046 57374 40102
rect 57430 40046 57498 40102
rect 57554 40046 57622 40102
rect 57678 40046 75250 40102
rect 75306 40046 75374 40102
rect 75430 40046 75498 40102
rect 75554 40046 75622 40102
rect 75678 40046 85238 40102
rect 85294 40046 85362 40102
rect 85418 40046 93250 40102
rect 93306 40046 93374 40102
rect 93430 40046 93498 40102
rect 93554 40046 93622 40102
rect 93678 40046 111250 40102
rect 111306 40046 111374 40102
rect 111430 40046 111498 40102
rect 111554 40046 111622 40102
rect 111678 40046 115958 40102
rect 116014 40046 116082 40102
rect 116138 40046 146678 40102
rect 146734 40046 146802 40102
rect 146858 40046 177398 40102
rect 177454 40046 177522 40102
rect 177578 40046 208118 40102
rect 208174 40046 208242 40102
rect 208298 40046 238838 40102
rect 238894 40046 238962 40102
rect 239018 40046 269558 40102
rect 269614 40046 269682 40102
rect 269738 40046 300278 40102
rect 300334 40046 300402 40102
rect 300458 40046 330998 40102
rect 331054 40046 331122 40102
rect 331178 40046 361718 40102
rect 361774 40046 361842 40102
rect 361898 40046 392438 40102
rect 392494 40046 392562 40102
rect 392618 40046 423158 40102
rect 423214 40046 423282 40102
rect 423338 40046 453878 40102
rect 453934 40046 454002 40102
rect 454058 40046 484598 40102
rect 484654 40046 484722 40102
rect 484778 40046 515318 40102
rect 515374 40046 515442 40102
rect 515498 40046 546038 40102
rect 546094 40046 546162 40102
rect 546218 40046 561250 40102
rect 561306 40046 561374 40102
rect 561430 40046 561498 40102
rect 561554 40046 561622 40102
rect 561678 40046 579250 40102
rect 579306 40046 579374 40102
rect 579430 40046 579498 40102
rect 579554 40046 579622 40102
rect 579678 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597980 40102
rect -1916 39978 597980 40046
rect -1916 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 3250 39978
rect 3306 39922 3374 39978
rect 3430 39922 3498 39978
rect 3554 39922 3622 39978
rect 3678 39922 21250 39978
rect 21306 39922 21374 39978
rect 21430 39922 21498 39978
rect 21554 39922 21622 39978
rect 21678 39922 39250 39978
rect 39306 39922 39374 39978
rect 39430 39922 39498 39978
rect 39554 39922 39622 39978
rect 39678 39922 54518 39978
rect 54574 39922 54642 39978
rect 54698 39922 57250 39978
rect 57306 39922 57374 39978
rect 57430 39922 57498 39978
rect 57554 39922 57622 39978
rect 57678 39922 75250 39978
rect 75306 39922 75374 39978
rect 75430 39922 75498 39978
rect 75554 39922 75622 39978
rect 75678 39922 85238 39978
rect 85294 39922 85362 39978
rect 85418 39922 93250 39978
rect 93306 39922 93374 39978
rect 93430 39922 93498 39978
rect 93554 39922 93622 39978
rect 93678 39922 111250 39978
rect 111306 39922 111374 39978
rect 111430 39922 111498 39978
rect 111554 39922 111622 39978
rect 111678 39922 115958 39978
rect 116014 39922 116082 39978
rect 116138 39922 146678 39978
rect 146734 39922 146802 39978
rect 146858 39922 177398 39978
rect 177454 39922 177522 39978
rect 177578 39922 208118 39978
rect 208174 39922 208242 39978
rect 208298 39922 238838 39978
rect 238894 39922 238962 39978
rect 239018 39922 269558 39978
rect 269614 39922 269682 39978
rect 269738 39922 300278 39978
rect 300334 39922 300402 39978
rect 300458 39922 330998 39978
rect 331054 39922 331122 39978
rect 331178 39922 361718 39978
rect 361774 39922 361842 39978
rect 361898 39922 392438 39978
rect 392494 39922 392562 39978
rect 392618 39922 423158 39978
rect 423214 39922 423282 39978
rect 423338 39922 453878 39978
rect 453934 39922 454002 39978
rect 454058 39922 484598 39978
rect 484654 39922 484722 39978
rect 484778 39922 515318 39978
rect 515374 39922 515442 39978
rect 515498 39922 546038 39978
rect 546094 39922 546162 39978
rect 546218 39922 561250 39978
rect 561306 39922 561374 39978
rect 561430 39922 561498 39978
rect 561554 39922 561622 39978
rect 561678 39922 579250 39978
rect 579306 39922 579374 39978
rect 579430 39922 579498 39978
rect 579554 39922 579622 39978
rect 579678 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597980 39978
rect -1916 39826 597980 39922
rect -1916 28350 597980 28446
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 6970 28350
rect 7026 28294 7094 28350
rect 7150 28294 7218 28350
rect 7274 28294 7342 28350
rect 7398 28294 24970 28350
rect 25026 28294 25094 28350
rect 25150 28294 25218 28350
rect 25274 28294 25342 28350
rect 25398 28294 42970 28350
rect 43026 28294 43094 28350
rect 43150 28294 43218 28350
rect 43274 28294 43342 28350
rect 43398 28294 60970 28350
rect 61026 28294 61094 28350
rect 61150 28294 61218 28350
rect 61274 28294 61342 28350
rect 61398 28294 78970 28350
rect 79026 28294 79094 28350
rect 79150 28294 79218 28350
rect 79274 28294 79342 28350
rect 79398 28294 96970 28350
rect 97026 28294 97094 28350
rect 97150 28294 97218 28350
rect 97274 28294 97342 28350
rect 97398 28294 114970 28350
rect 115026 28294 115094 28350
rect 115150 28294 115218 28350
rect 115274 28294 115342 28350
rect 115398 28294 132970 28350
rect 133026 28294 133094 28350
rect 133150 28294 133218 28350
rect 133274 28294 133342 28350
rect 133398 28294 150970 28350
rect 151026 28294 151094 28350
rect 151150 28294 151218 28350
rect 151274 28294 151342 28350
rect 151398 28294 168970 28350
rect 169026 28294 169094 28350
rect 169150 28294 169218 28350
rect 169274 28294 169342 28350
rect 169398 28294 186970 28350
rect 187026 28294 187094 28350
rect 187150 28294 187218 28350
rect 187274 28294 187342 28350
rect 187398 28294 204970 28350
rect 205026 28294 205094 28350
rect 205150 28294 205218 28350
rect 205274 28294 205342 28350
rect 205398 28294 222970 28350
rect 223026 28294 223094 28350
rect 223150 28294 223218 28350
rect 223274 28294 223342 28350
rect 223398 28294 240970 28350
rect 241026 28294 241094 28350
rect 241150 28294 241218 28350
rect 241274 28294 241342 28350
rect 241398 28294 258970 28350
rect 259026 28294 259094 28350
rect 259150 28294 259218 28350
rect 259274 28294 259342 28350
rect 259398 28294 276970 28350
rect 277026 28294 277094 28350
rect 277150 28294 277218 28350
rect 277274 28294 277342 28350
rect 277398 28294 294970 28350
rect 295026 28294 295094 28350
rect 295150 28294 295218 28350
rect 295274 28294 295342 28350
rect 295398 28294 312970 28350
rect 313026 28294 313094 28350
rect 313150 28294 313218 28350
rect 313274 28294 313342 28350
rect 313398 28294 330970 28350
rect 331026 28294 331094 28350
rect 331150 28294 331218 28350
rect 331274 28294 331342 28350
rect 331398 28294 348970 28350
rect 349026 28294 349094 28350
rect 349150 28294 349218 28350
rect 349274 28294 349342 28350
rect 349398 28294 366970 28350
rect 367026 28294 367094 28350
rect 367150 28294 367218 28350
rect 367274 28294 367342 28350
rect 367398 28294 384970 28350
rect 385026 28294 385094 28350
rect 385150 28294 385218 28350
rect 385274 28294 385342 28350
rect 385398 28294 402970 28350
rect 403026 28294 403094 28350
rect 403150 28294 403218 28350
rect 403274 28294 403342 28350
rect 403398 28294 420970 28350
rect 421026 28294 421094 28350
rect 421150 28294 421218 28350
rect 421274 28294 421342 28350
rect 421398 28294 438970 28350
rect 439026 28294 439094 28350
rect 439150 28294 439218 28350
rect 439274 28294 439342 28350
rect 439398 28294 456970 28350
rect 457026 28294 457094 28350
rect 457150 28294 457218 28350
rect 457274 28294 457342 28350
rect 457398 28294 474970 28350
rect 475026 28294 475094 28350
rect 475150 28294 475218 28350
rect 475274 28294 475342 28350
rect 475398 28294 492970 28350
rect 493026 28294 493094 28350
rect 493150 28294 493218 28350
rect 493274 28294 493342 28350
rect 493398 28294 510970 28350
rect 511026 28294 511094 28350
rect 511150 28294 511218 28350
rect 511274 28294 511342 28350
rect 511398 28294 528970 28350
rect 529026 28294 529094 28350
rect 529150 28294 529218 28350
rect 529274 28294 529342 28350
rect 529398 28294 546970 28350
rect 547026 28294 547094 28350
rect 547150 28294 547218 28350
rect 547274 28294 547342 28350
rect 547398 28294 564970 28350
rect 565026 28294 565094 28350
rect 565150 28294 565218 28350
rect 565274 28294 565342 28350
rect 565398 28294 582970 28350
rect 583026 28294 583094 28350
rect 583150 28294 583218 28350
rect 583274 28294 583342 28350
rect 583398 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect -1916 28226 597980 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 6970 28226
rect 7026 28170 7094 28226
rect 7150 28170 7218 28226
rect 7274 28170 7342 28226
rect 7398 28170 24970 28226
rect 25026 28170 25094 28226
rect 25150 28170 25218 28226
rect 25274 28170 25342 28226
rect 25398 28170 42970 28226
rect 43026 28170 43094 28226
rect 43150 28170 43218 28226
rect 43274 28170 43342 28226
rect 43398 28170 60970 28226
rect 61026 28170 61094 28226
rect 61150 28170 61218 28226
rect 61274 28170 61342 28226
rect 61398 28170 78970 28226
rect 79026 28170 79094 28226
rect 79150 28170 79218 28226
rect 79274 28170 79342 28226
rect 79398 28170 96970 28226
rect 97026 28170 97094 28226
rect 97150 28170 97218 28226
rect 97274 28170 97342 28226
rect 97398 28170 114970 28226
rect 115026 28170 115094 28226
rect 115150 28170 115218 28226
rect 115274 28170 115342 28226
rect 115398 28170 132970 28226
rect 133026 28170 133094 28226
rect 133150 28170 133218 28226
rect 133274 28170 133342 28226
rect 133398 28170 150970 28226
rect 151026 28170 151094 28226
rect 151150 28170 151218 28226
rect 151274 28170 151342 28226
rect 151398 28170 168970 28226
rect 169026 28170 169094 28226
rect 169150 28170 169218 28226
rect 169274 28170 169342 28226
rect 169398 28170 186970 28226
rect 187026 28170 187094 28226
rect 187150 28170 187218 28226
rect 187274 28170 187342 28226
rect 187398 28170 204970 28226
rect 205026 28170 205094 28226
rect 205150 28170 205218 28226
rect 205274 28170 205342 28226
rect 205398 28170 222970 28226
rect 223026 28170 223094 28226
rect 223150 28170 223218 28226
rect 223274 28170 223342 28226
rect 223398 28170 240970 28226
rect 241026 28170 241094 28226
rect 241150 28170 241218 28226
rect 241274 28170 241342 28226
rect 241398 28170 258970 28226
rect 259026 28170 259094 28226
rect 259150 28170 259218 28226
rect 259274 28170 259342 28226
rect 259398 28170 276970 28226
rect 277026 28170 277094 28226
rect 277150 28170 277218 28226
rect 277274 28170 277342 28226
rect 277398 28170 294970 28226
rect 295026 28170 295094 28226
rect 295150 28170 295218 28226
rect 295274 28170 295342 28226
rect 295398 28170 312970 28226
rect 313026 28170 313094 28226
rect 313150 28170 313218 28226
rect 313274 28170 313342 28226
rect 313398 28170 330970 28226
rect 331026 28170 331094 28226
rect 331150 28170 331218 28226
rect 331274 28170 331342 28226
rect 331398 28170 348970 28226
rect 349026 28170 349094 28226
rect 349150 28170 349218 28226
rect 349274 28170 349342 28226
rect 349398 28170 366970 28226
rect 367026 28170 367094 28226
rect 367150 28170 367218 28226
rect 367274 28170 367342 28226
rect 367398 28170 384970 28226
rect 385026 28170 385094 28226
rect 385150 28170 385218 28226
rect 385274 28170 385342 28226
rect 385398 28170 402970 28226
rect 403026 28170 403094 28226
rect 403150 28170 403218 28226
rect 403274 28170 403342 28226
rect 403398 28170 420970 28226
rect 421026 28170 421094 28226
rect 421150 28170 421218 28226
rect 421274 28170 421342 28226
rect 421398 28170 438970 28226
rect 439026 28170 439094 28226
rect 439150 28170 439218 28226
rect 439274 28170 439342 28226
rect 439398 28170 456970 28226
rect 457026 28170 457094 28226
rect 457150 28170 457218 28226
rect 457274 28170 457342 28226
rect 457398 28170 474970 28226
rect 475026 28170 475094 28226
rect 475150 28170 475218 28226
rect 475274 28170 475342 28226
rect 475398 28170 492970 28226
rect 493026 28170 493094 28226
rect 493150 28170 493218 28226
rect 493274 28170 493342 28226
rect 493398 28170 510970 28226
rect 511026 28170 511094 28226
rect 511150 28170 511218 28226
rect 511274 28170 511342 28226
rect 511398 28170 528970 28226
rect 529026 28170 529094 28226
rect 529150 28170 529218 28226
rect 529274 28170 529342 28226
rect 529398 28170 546970 28226
rect 547026 28170 547094 28226
rect 547150 28170 547218 28226
rect 547274 28170 547342 28226
rect 547398 28170 564970 28226
rect 565026 28170 565094 28226
rect 565150 28170 565218 28226
rect 565274 28170 565342 28226
rect 565398 28170 582970 28226
rect 583026 28170 583094 28226
rect 583150 28170 583218 28226
rect 583274 28170 583342 28226
rect 583398 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect -1916 28102 597980 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 6970 28102
rect 7026 28046 7094 28102
rect 7150 28046 7218 28102
rect 7274 28046 7342 28102
rect 7398 28046 24970 28102
rect 25026 28046 25094 28102
rect 25150 28046 25218 28102
rect 25274 28046 25342 28102
rect 25398 28046 42970 28102
rect 43026 28046 43094 28102
rect 43150 28046 43218 28102
rect 43274 28046 43342 28102
rect 43398 28046 60970 28102
rect 61026 28046 61094 28102
rect 61150 28046 61218 28102
rect 61274 28046 61342 28102
rect 61398 28046 78970 28102
rect 79026 28046 79094 28102
rect 79150 28046 79218 28102
rect 79274 28046 79342 28102
rect 79398 28046 96970 28102
rect 97026 28046 97094 28102
rect 97150 28046 97218 28102
rect 97274 28046 97342 28102
rect 97398 28046 114970 28102
rect 115026 28046 115094 28102
rect 115150 28046 115218 28102
rect 115274 28046 115342 28102
rect 115398 28046 132970 28102
rect 133026 28046 133094 28102
rect 133150 28046 133218 28102
rect 133274 28046 133342 28102
rect 133398 28046 150970 28102
rect 151026 28046 151094 28102
rect 151150 28046 151218 28102
rect 151274 28046 151342 28102
rect 151398 28046 168970 28102
rect 169026 28046 169094 28102
rect 169150 28046 169218 28102
rect 169274 28046 169342 28102
rect 169398 28046 186970 28102
rect 187026 28046 187094 28102
rect 187150 28046 187218 28102
rect 187274 28046 187342 28102
rect 187398 28046 204970 28102
rect 205026 28046 205094 28102
rect 205150 28046 205218 28102
rect 205274 28046 205342 28102
rect 205398 28046 222970 28102
rect 223026 28046 223094 28102
rect 223150 28046 223218 28102
rect 223274 28046 223342 28102
rect 223398 28046 240970 28102
rect 241026 28046 241094 28102
rect 241150 28046 241218 28102
rect 241274 28046 241342 28102
rect 241398 28046 258970 28102
rect 259026 28046 259094 28102
rect 259150 28046 259218 28102
rect 259274 28046 259342 28102
rect 259398 28046 276970 28102
rect 277026 28046 277094 28102
rect 277150 28046 277218 28102
rect 277274 28046 277342 28102
rect 277398 28046 294970 28102
rect 295026 28046 295094 28102
rect 295150 28046 295218 28102
rect 295274 28046 295342 28102
rect 295398 28046 312970 28102
rect 313026 28046 313094 28102
rect 313150 28046 313218 28102
rect 313274 28046 313342 28102
rect 313398 28046 330970 28102
rect 331026 28046 331094 28102
rect 331150 28046 331218 28102
rect 331274 28046 331342 28102
rect 331398 28046 348970 28102
rect 349026 28046 349094 28102
rect 349150 28046 349218 28102
rect 349274 28046 349342 28102
rect 349398 28046 366970 28102
rect 367026 28046 367094 28102
rect 367150 28046 367218 28102
rect 367274 28046 367342 28102
rect 367398 28046 384970 28102
rect 385026 28046 385094 28102
rect 385150 28046 385218 28102
rect 385274 28046 385342 28102
rect 385398 28046 402970 28102
rect 403026 28046 403094 28102
rect 403150 28046 403218 28102
rect 403274 28046 403342 28102
rect 403398 28046 420970 28102
rect 421026 28046 421094 28102
rect 421150 28046 421218 28102
rect 421274 28046 421342 28102
rect 421398 28046 438970 28102
rect 439026 28046 439094 28102
rect 439150 28046 439218 28102
rect 439274 28046 439342 28102
rect 439398 28046 456970 28102
rect 457026 28046 457094 28102
rect 457150 28046 457218 28102
rect 457274 28046 457342 28102
rect 457398 28046 474970 28102
rect 475026 28046 475094 28102
rect 475150 28046 475218 28102
rect 475274 28046 475342 28102
rect 475398 28046 492970 28102
rect 493026 28046 493094 28102
rect 493150 28046 493218 28102
rect 493274 28046 493342 28102
rect 493398 28046 510970 28102
rect 511026 28046 511094 28102
rect 511150 28046 511218 28102
rect 511274 28046 511342 28102
rect 511398 28046 528970 28102
rect 529026 28046 529094 28102
rect 529150 28046 529218 28102
rect 529274 28046 529342 28102
rect 529398 28046 546970 28102
rect 547026 28046 547094 28102
rect 547150 28046 547218 28102
rect 547274 28046 547342 28102
rect 547398 28046 564970 28102
rect 565026 28046 565094 28102
rect 565150 28046 565218 28102
rect 565274 28046 565342 28102
rect 565398 28046 582970 28102
rect 583026 28046 583094 28102
rect 583150 28046 583218 28102
rect 583274 28046 583342 28102
rect 583398 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect -1916 27978 597980 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 6970 27978
rect 7026 27922 7094 27978
rect 7150 27922 7218 27978
rect 7274 27922 7342 27978
rect 7398 27922 24970 27978
rect 25026 27922 25094 27978
rect 25150 27922 25218 27978
rect 25274 27922 25342 27978
rect 25398 27922 42970 27978
rect 43026 27922 43094 27978
rect 43150 27922 43218 27978
rect 43274 27922 43342 27978
rect 43398 27922 60970 27978
rect 61026 27922 61094 27978
rect 61150 27922 61218 27978
rect 61274 27922 61342 27978
rect 61398 27922 78970 27978
rect 79026 27922 79094 27978
rect 79150 27922 79218 27978
rect 79274 27922 79342 27978
rect 79398 27922 96970 27978
rect 97026 27922 97094 27978
rect 97150 27922 97218 27978
rect 97274 27922 97342 27978
rect 97398 27922 114970 27978
rect 115026 27922 115094 27978
rect 115150 27922 115218 27978
rect 115274 27922 115342 27978
rect 115398 27922 132970 27978
rect 133026 27922 133094 27978
rect 133150 27922 133218 27978
rect 133274 27922 133342 27978
rect 133398 27922 150970 27978
rect 151026 27922 151094 27978
rect 151150 27922 151218 27978
rect 151274 27922 151342 27978
rect 151398 27922 168970 27978
rect 169026 27922 169094 27978
rect 169150 27922 169218 27978
rect 169274 27922 169342 27978
rect 169398 27922 186970 27978
rect 187026 27922 187094 27978
rect 187150 27922 187218 27978
rect 187274 27922 187342 27978
rect 187398 27922 204970 27978
rect 205026 27922 205094 27978
rect 205150 27922 205218 27978
rect 205274 27922 205342 27978
rect 205398 27922 222970 27978
rect 223026 27922 223094 27978
rect 223150 27922 223218 27978
rect 223274 27922 223342 27978
rect 223398 27922 240970 27978
rect 241026 27922 241094 27978
rect 241150 27922 241218 27978
rect 241274 27922 241342 27978
rect 241398 27922 258970 27978
rect 259026 27922 259094 27978
rect 259150 27922 259218 27978
rect 259274 27922 259342 27978
rect 259398 27922 276970 27978
rect 277026 27922 277094 27978
rect 277150 27922 277218 27978
rect 277274 27922 277342 27978
rect 277398 27922 294970 27978
rect 295026 27922 295094 27978
rect 295150 27922 295218 27978
rect 295274 27922 295342 27978
rect 295398 27922 312970 27978
rect 313026 27922 313094 27978
rect 313150 27922 313218 27978
rect 313274 27922 313342 27978
rect 313398 27922 330970 27978
rect 331026 27922 331094 27978
rect 331150 27922 331218 27978
rect 331274 27922 331342 27978
rect 331398 27922 348970 27978
rect 349026 27922 349094 27978
rect 349150 27922 349218 27978
rect 349274 27922 349342 27978
rect 349398 27922 366970 27978
rect 367026 27922 367094 27978
rect 367150 27922 367218 27978
rect 367274 27922 367342 27978
rect 367398 27922 384970 27978
rect 385026 27922 385094 27978
rect 385150 27922 385218 27978
rect 385274 27922 385342 27978
rect 385398 27922 402970 27978
rect 403026 27922 403094 27978
rect 403150 27922 403218 27978
rect 403274 27922 403342 27978
rect 403398 27922 420970 27978
rect 421026 27922 421094 27978
rect 421150 27922 421218 27978
rect 421274 27922 421342 27978
rect 421398 27922 438970 27978
rect 439026 27922 439094 27978
rect 439150 27922 439218 27978
rect 439274 27922 439342 27978
rect 439398 27922 456970 27978
rect 457026 27922 457094 27978
rect 457150 27922 457218 27978
rect 457274 27922 457342 27978
rect 457398 27922 474970 27978
rect 475026 27922 475094 27978
rect 475150 27922 475218 27978
rect 475274 27922 475342 27978
rect 475398 27922 492970 27978
rect 493026 27922 493094 27978
rect 493150 27922 493218 27978
rect 493274 27922 493342 27978
rect 493398 27922 510970 27978
rect 511026 27922 511094 27978
rect 511150 27922 511218 27978
rect 511274 27922 511342 27978
rect 511398 27922 528970 27978
rect 529026 27922 529094 27978
rect 529150 27922 529218 27978
rect 529274 27922 529342 27978
rect 529398 27922 546970 27978
rect 547026 27922 547094 27978
rect 547150 27922 547218 27978
rect 547274 27922 547342 27978
rect 547398 27922 564970 27978
rect 565026 27922 565094 27978
rect 565150 27922 565218 27978
rect 565274 27922 565342 27978
rect 565398 27922 582970 27978
rect 583026 27922 583094 27978
rect 583150 27922 583218 27978
rect 583274 27922 583342 27978
rect 583398 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect -1916 27826 597980 27922
rect -1916 22350 597980 22446
rect -1916 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 3250 22350
rect 3306 22294 3374 22350
rect 3430 22294 3498 22350
rect 3554 22294 3622 22350
rect 3678 22294 21250 22350
rect 21306 22294 21374 22350
rect 21430 22294 21498 22350
rect 21554 22294 21622 22350
rect 21678 22294 39250 22350
rect 39306 22294 39374 22350
rect 39430 22294 39498 22350
rect 39554 22294 39622 22350
rect 39678 22294 57250 22350
rect 57306 22294 57374 22350
rect 57430 22294 57498 22350
rect 57554 22294 57622 22350
rect 57678 22294 75250 22350
rect 75306 22294 75374 22350
rect 75430 22294 75498 22350
rect 75554 22294 75622 22350
rect 75678 22294 93250 22350
rect 93306 22294 93374 22350
rect 93430 22294 93498 22350
rect 93554 22294 93622 22350
rect 93678 22294 111250 22350
rect 111306 22294 111374 22350
rect 111430 22294 111498 22350
rect 111554 22294 111622 22350
rect 111678 22294 129250 22350
rect 129306 22294 129374 22350
rect 129430 22294 129498 22350
rect 129554 22294 129622 22350
rect 129678 22294 147250 22350
rect 147306 22294 147374 22350
rect 147430 22294 147498 22350
rect 147554 22294 147622 22350
rect 147678 22294 165250 22350
rect 165306 22294 165374 22350
rect 165430 22294 165498 22350
rect 165554 22294 165622 22350
rect 165678 22294 183250 22350
rect 183306 22294 183374 22350
rect 183430 22294 183498 22350
rect 183554 22294 183622 22350
rect 183678 22294 201250 22350
rect 201306 22294 201374 22350
rect 201430 22294 201498 22350
rect 201554 22294 201622 22350
rect 201678 22294 219250 22350
rect 219306 22294 219374 22350
rect 219430 22294 219498 22350
rect 219554 22294 219622 22350
rect 219678 22294 237250 22350
rect 237306 22294 237374 22350
rect 237430 22294 237498 22350
rect 237554 22294 237622 22350
rect 237678 22294 255250 22350
rect 255306 22294 255374 22350
rect 255430 22294 255498 22350
rect 255554 22294 255622 22350
rect 255678 22294 273250 22350
rect 273306 22294 273374 22350
rect 273430 22294 273498 22350
rect 273554 22294 273622 22350
rect 273678 22294 291250 22350
rect 291306 22294 291374 22350
rect 291430 22294 291498 22350
rect 291554 22294 291622 22350
rect 291678 22294 309250 22350
rect 309306 22294 309374 22350
rect 309430 22294 309498 22350
rect 309554 22294 309622 22350
rect 309678 22294 327250 22350
rect 327306 22294 327374 22350
rect 327430 22294 327498 22350
rect 327554 22294 327622 22350
rect 327678 22294 345250 22350
rect 345306 22294 345374 22350
rect 345430 22294 345498 22350
rect 345554 22294 345622 22350
rect 345678 22294 363250 22350
rect 363306 22294 363374 22350
rect 363430 22294 363498 22350
rect 363554 22294 363622 22350
rect 363678 22294 381250 22350
rect 381306 22294 381374 22350
rect 381430 22294 381498 22350
rect 381554 22294 381622 22350
rect 381678 22294 399250 22350
rect 399306 22294 399374 22350
rect 399430 22294 399498 22350
rect 399554 22294 399622 22350
rect 399678 22294 417250 22350
rect 417306 22294 417374 22350
rect 417430 22294 417498 22350
rect 417554 22294 417622 22350
rect 417678 22294 435250 22350
rect 435306 22294 435374 22350
rect 435430 22294 435498 22350
rect 435554 22294 435622 22350
rect 435678 22294 453250 22350
rect 453306 22294 453374 22350
rect 453430 22294 453498 22350
rect 453554 22294 453622 22350
rect 453678 22294 471250 22350
rect 471306 22294 471374 22350
rect 471430 22294 471498 22350
rect 471554 22294 471622 22350
rect 471678 22294 489250 22350
rect 489306 22294 489374 22350
rect 489430 22294 489498 22350
rect 489554 22294 489622 22350
rect 489678 22294 507250 22350
rect 507306 22294 507374 22350
rect 507430 22294 507498 22350
rect 507554 22294 507622 22350
rect 507678 22294 525250 22350
rect 525306 22294 525374 22350
rect 525430 22294 525498 22350
rect 525554 22294 525622 22350
rect 525678 22294 543250 22350
rect 543306 22294 543374 22350
rect 543430 22294 543498 22350
rect 543554 22294 543622 22350
rect 543678 22294 561250 22350
rect 561306 22294 561374 22350
rect 561430 22294 561498 22350
rect 561554 22294 561622 22350
rect 561678 22294 579250 22350
rect 579306 22294 579374 22350
rect 579430 22294 579498 22350
rect 579554 22294 579622 22350
rect 579678 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597980 22350
rect -1916 22226 597980 22294
rect -1916 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 3250 22226
rect 3306 22170 3374 22226
rect 3430 22170 3498 22226
rect 3554 22170 3622 22226
rect 3678 22170 21250 22226
rect 21306 22170 21374 22226
rect 21430 22170 21498 22226
rect 21554 22170 21622 22226
rect 21678 22170 39250 22226
rect 39306 22170 39374 22226
rect 39430 22170 39498 22226
rect 39554 22170 39622 22226
rect 39678 22170 57250 22226
rect 57306 22170 57374 22226
rect 57430 22170 57498 22226
rect 57554 22170 57622 22226
rect 57678 22170 75250 22226
rect 75306 22170 75374 22226
rect 75430 22170 75498 22226
rect 75554 22170 75622 22226
rect 75678 22170 93250 22226
rect 93306 22170 93374 22226
rect 93430 22170 93498 22226
rect 93554 22170 93622 22226
rect 93678 22170 111250 22226
rect 111306 22170 111374 22226
rect 111430 22170 111498 22226
rect 111554 22170 111622 22226
rect 111678 22170 129250 22226
rect 129306 22170 129374 22226
rect 129430 22170 129498 22226
rect 129554 22170 129622 22226
rect 129678 22170 147250 22226
rect 147306 22170 147374 22226
rect 147430 22170 147498 22226
rect 147554 22170 147622 22226
rect 147678 22170 165250 22226
rect 165306 22170 165374 22226
rect 165430 22170 165498 22226
rect 165554 22170 165622 22226
rect 165678 22170 183250 22226
rect 183306 22170 183374 22226
rect 183430 22170 183498 22226
rect 183554 22170 183622 22226
rect 183678 22170 201250 22226
rect 201306 22170 201374 22226
rect 201430 22170 201498 22226
rect 201554 22170 201622 22226
rect 201678 22170 219250 22226
rect 219306 22170 219374 22226
rect 219430 22170 219498 22226
rect 219554 22170 219622 22226
rect 219678 22170 237250 22226
rect 237306 22170 237374 22226
rect 237430 22170 237498 22226
rect 237554 22170 237622 22226
rect 237678 22170 255250 22226
rect 255306 22170 255374 22226
rect 255430 22170 255498 22226
rect 255554 22170 255622 22226
rect 255678 22170 273250 22226
rect 273306 22170 273374 22226
rect 273430 22170 273498 22226
rect 273554 22170 273622 22226
rect 273678 22170 291250 22226
rect 291306 22170 291374 22226
rect 291430 22170 291498 22226
rect 291554 22170 291622 22226
rect 291678 22170 309250 22226
rect 309306 22170 309374 22226
rect 309430 22170 309498 22226
rect 309554 22170 309622 22226
rect 309678 22170 327250 22226
rect 327306 22170 327374 22226
rect 327430 22170 327498 22226
rect 327554 22170 327622 22226
rect 327678 22170 345250 22226
rect 345306 22170 345374 22226
rect 345430 22170 345498 22226
rect 345554 22170 345622 22226
rect 345678 22170 363250 22226
rect 363306 22170 363374 22226
rect 363430 22170 363498 22226
rect 363554 22170 363622 22226
rect 363678 22170 381250 22226
rect 381306 22170 381374 22226
rect 381430 22170 381498 22226
rect 381554 22170 381622 22226
rect 381678 22170 399250 22226
rect 399306 22170 399374 22226
rect 399430 22170 399498 22226
rect 399554 22170 399622 22226
rect 399678 22170 417250 22226
rect 417306 22170 417374 22226
rect 417430 22170 417498 22226
rect 417554 22170 417622 22226
rect 417678 22170 435250 22226
rect 435306 22170 435374 22226
rect 435430 22170 435498 22226
rect 435554 22170 435622 22226
rect 435678 22170 453250 22226
rect 453306 22170 453374 22226
rect 453430 22170 453498 22226
rect 453554 22170 453622 22226
rect 453678 22170 471250 22226
rect 471306 22170 471374 22226
rect 471430 22170 471498 22226
rect 471554 22170 471622 22226
rect 471678 22170 489250 22226
rect 489306 22170 489374 22226
rect 489430 22170 489498 22226
rect 489554 22170 489622 22226
rect 489678 22170 507250 22226
rect 507306 22170 507374 22226
rect 507430 22170 507498 22226
rect 507554 22170 507622 22226
rect 507678 22170 525250 22226
rect 525306 22170 525374 22226
rect 525430 22170 525498 22226
rect 525554 22170 525622 22226
rect 525678 22170 543250 22226
rect 543306 22170 543374 22226
rect 543430 22170 543498 22226
rect 543554 22170 543622 22226
rect 543678 22170 561250 22226
rect 561306 22170 561374 22226
rect 561430 22170 561498 22226
rect 561554 22170 561622 22226
rect 561678 22170 579250 22226
rect 579306 22170 579374 22226
rect 579430 22170 579498 22226
rect 579554 22170 579622 22226
rect 579678 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597980 22226
rect -1916 22102 597980 22170
rect -1916 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 3250 22102
rect 3306 22046 3374 22102
rect 3430 22046 3498 22102
rect 3554 22046 3622 22102
rect 3678 22046 21250 22102
rect 21306 22046 21374 22102
rect 21430 22046 21498 22102
rect 21554 22046 21622 22102
rect 21678 22046 39250 22102
rect 39306 22046 39374 22102
rect 39430 22046 39498 22102
rect 39554 22046 39622 22102
rect 39678 22046 57250 22102
rect 57306 22046 57374 22102
rect 57430 22046 57498 22102
rect 57554 22046 57622 22102
rect 57678 22046 75250 22102
rect 75306 22046 75374 22102
rect 75430 22046 75498 22102
rect 75554 22046 75622 22102
rect 75678 22046 93250 22102
rect 93306 22046 93374 22102
rect 93430 22046 93498 22102
rect 93554 22046 93622 22102
rect 93678 22046 111250 22102
rect 111306 22046 111374 22102
rect 111430 22046 111498 22102
rect 111554 22046 111622 22102
rect 111678 22046 129250 22102
rect 129306 22046 129374 22102
rect 129430 22046 129498 22102
rect 129554 22046 129622 22102
rect 129678 22046 147250 22102
rect 147306 22046 147374 22102
rect 147430 22046 147498 22102
rect 147554 22046 147622 22102
rect 147678 22046 165250 22102
rect 165306 22046 165374 22102
rect 165430 22046 165498 22102
rect 165554 22046 165622 22102
rect 165678 22046 183250 22102
rect 183306 22046 183374 22102
rect 183430 22046 183498 22102
rect 183554 22046 183622 22102
rect 183678 22046 201250 22102
rect 201306 22046 201374 22102
rect 201430 22046 201498 22102
rect 201554 22046 201622 22102
rect 201678 22046 219250 22102
rect 219306 22046 219374 22102
rect 219430 22046 219498 22102
rect 219554 22046 219622 22102
rect 219678 22046 237250 22102
rect 237306 22046 237374 22102
rect 237430 22046 237498 22102
rect 237554 22046 237622 22102
rect 237678 22046 255250 22102
rect 255306 22046 255374 22102
rect 255430 22046 255498 22102
rect 255554 22046 255622 22102
rect 255678 22046 273250 22102
rect 273306 22046 273374 22102
rect 273430 22046 273498 22102
rect 273554 22046 273622 22102
rect 273678 22046 291250 22102
rect 291306 22046 291374 22102
rect 291430 22046 291498 22102
rect 291554 22046 291622 22102
rect 291678 22046 309250 22102
rect 309306 22046 309374 22102
rect 309430 22046 309498 22102
rect 309554 22046 309622 22102
rect 309678 22046 327250 22102
rect 327306 22046 327374 22102
rect 327430 22046 327498 22102
rect 327554 22046 327622 22102
rect 327678 22046 345250 22102
rect 345306 22046 345374 22102
rect 345430 22046 345498 22102
rect 345554 22046 345622 22102
rect 345678 22046 363250 22102
rect 363306 22046 363374 22102
rect 363430 22046 363498 22102
rect 363554 22046 363622 22102
rect 363678 22046 381250 22102
rect 381306 22046 381374 22102
rect 381430 22046 381498 22102
rect 381554 22046 381622 22102
rect 381678 22046 399250 22102
rect 399306 22046 399374 22102
rect 399430 22046 399498 22102
rect 399554 22046 399622 22102
rect 399678 22046 417250 22102
rect 417306 22046 417374 22102
rect 417430 22046 417498 22102
rect 417554 22046 417622 22102
rect 417678 22046 435250 22102
rect 435306 22046 435374 22102
rect 435430 22046 435498 22102
rect 435554 22046 435622 22102
rect 435678 22046 453250 22102
rect 453306 22046 453374 22102
rect 453430 22046 453498 22102
rect 453554 22046 453622 22102
rect 453678 22046 471250 22102
rect 471306 22046 471374 22102
rect 471430 22046 471498 22102
rect 471554 22046 471622 22102
rect 471678 22046 489250 22102
rect 489306 22046 489374 22102
rect 489430 22046 489498 22102
rect 489554 22046 489622 22102
rect 489678 22046 507250 22102
rect 507306 22046 507374 22102
rect 507430 22046 507498 22102
rect 507554 22046 507622 22102
rect 507678 22046 525250 22102
rect 525306 22046 525374 22102
rect 525430 22046 525498 22102
rect 525554 22046 525622 22102
rect 525678 22046 543250 22102
rect 543306 22046 543374 22102
rect 543430 22046 543498 22102
rect 543554 22046 543622 22102
rect 543678 22046 561250 22102
rect 561306 22046 561374 22102
rect 561430 22046 561498 22102
rect 561554 22046 561622 22102
rect 561678 22046 579250 22102
rect 579306 22046 579374 22102
rect 579430 22046 579498 22102
rect 579554 22046 579622 22102
rect 579678 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597980 22102
rect -1916 21978 597980 22046
rect -1916 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 3250 21978
rect 3306 21922 3374 21978
rect 3430 21922 3498 21978
rect 3554 21922 3622 21978
rect 3678 21922 21250 21978
rect 21306 21922 21374 21978
rect 21430 21922 21498 21978
rect 21554 21922 21622 21978
rect 21678 21922 39250 21978
rect 39306 21922 39374 21978
rect 39430 21922 39498 21978
rect 39554 21922 39622 21978
rect 39678 21922 57250 21978
rect 57306 21922 57374 21978
rect 57430 21922 57498 21978
rect 57554 21922 57622 21978
rect 57678 21922 75250 21978
rect 75306 21922 75374 21978
rect 75430 21922 75498 21978
rect 75554 21922 75622 21978
rect 75678 21922 93250 21978
rect 93306 21922 93374 21978
rect 93430 21922 93498 21978
rect 93554 21922 93622 21978
rect 93678 21922 111250 21978
rect 111306 21922 111374 21978
rect 111430 21922 111498 21978
rect 111554 21922 111622 21978
rect 111678 21922 129250 21978
rect 129306 21922 129374 21978
rect 129430 21922 129498 21978
rect 129554 21922 129622 21978
rect 129678 21922 147250 21978
rect 147306 21922 147374 21978
rect 147430 21922 147498 21978
rect 147554 21922 147622 21978
rect 147678 21922 165250 21978
rect 165306 21922 165374 21978
rect 165430 21922 165498 21978
rect 165554 21922 165622 21978
rect 165678 21922 183250 21978
rect 183306 21922 183374 21978
rect 183430 21922 183498 21978
rect 183554 21922 183622 21978
rect 183678 21922 201250 21978
rect 201306 21922 201374 21978
rect 201430 21922 201498 21978
rect 201554 21922 201622 21978
rect 201678 21922 219250 21978
rect 219306 21922 219374 21978
rect 219430 21922 219498 21978
rect 219554 21922 219622 21978
rect 219678 21922 237250 21978
rect 237306 21922 237374 21978
rect 237430 21922 237498 21978
rect 237554 21922 237622 21978
rect 237678 21922 255250 21978
rect 255306 21922 255374 21978
rect 255430 21922 255498 21978
rect 255554 21922 255622 21978
rect 255678 21922 273250 21978
rect 273306 21922 273374 21978
rect 273430 21922 273498 21978
rect 273554 21922 273622 21978
rect 273678 21922 291250 21978
rect 291306 21922 291374 21978
rect 291430 21922 291498 21978
rect 291554 21922 291622 21978
rect 291678 21922 309250 21978
rect 309306 21922 309374 21978
rect 309430 21922 309498 21978
rect 309554 21922 309622 21978
rect 309678 21922 327250 21978
rect 327306 21922 327374 21978
rect 327430 21922 327498 21978
rect 327554 21922 327622 21978
rect 327678 21922 345250 21978
rect 345306 21922 345374 21978
rect 345430 21922 345498 21978
rect 345554 21922 345622 21978
rect 345678 21922 363250 21978
rect 363306 21922 363374 21978
rect 363430 21922 363498 21978
rect 363554 21922 363622 21978
rect 363678 21922 381250 21978
rect 381306 21922 381374 21978
rect 381430 21922 381498 21978
rect 381554 21922 381622 21978
rect 381678 21922 399250 21978
rect 399306 21922 399374 21978
rect 399430 21922 399498 21978
rect 399554 21922 399622 21978
rect 399678 21922 417250 21978
rect 417306 21922 417374 21978
rect 417430 21922 417498 21978
rect 417554 21922 417622 21978
rect 417678 21922 435250 21978
rect 435306 21922 435374 21978
rect 435430 21922 435498 21978
rect 435554 21922 435622 21978
rect 435678 21922 453250 21978
rect 453306 21922 453374 21978
rect 453430 21922 453498 21978
rect 453554 21922 453622 21978
rect 453678 21922 471250 21978
rect 471306 21922 471374 21978
rect 471430 21922 471498 21978
rect 471554 21922 471622 21978
rect 471678 21922 489250 21978
rect 489306 21922 489374 21978
rect 489430 21922 489498 21978
rect 489554 21922 489622 21978
rect 489678 21922 507250 21978
rect 507306 21922 507374 21978
rect 507430 21922 507498 21978
rect 507554 21922 507622 21978
rect 507678 21922 525250 21978
rect 525306 21922 525374 21978
rect 525430 21922 525498 21978
rect 525554 21922 525622 21978
rect 525678 21922 543250 21978
rect 543306 21922 543374 21978
rect 543430 21922 543498 21978
rect 543554 21922 543622 21978
rect 543678 21922 561250 21978
rect 561306 21922 561374 21978
rect 561430 21922 561498 21978
rect 561554 21922 561622 21978
rect 561678 21922 579250 21978
rect 579306 21922 579374 21978
rect 579430 21922 579498 21978
rect 579554 21922 579622 21978
rect 579678 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597980 21978
rect -1916 21826 597980 21922
rect -1916 10350 597980 10446
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 6970 10350
rect 7026 10294 7094 10350
rect 7150 10294 7218 10350
rect 7274 10294 7342 10350
rect 7398 10294 24970 10350
rect 25026 10294 25094 10350
rect 25150 10294 25218 10350
rect 25274 10294 25342 10350
rect 25398 10294 42970 10350
rect 43026 10294 43094 10350
rect 43150 10294 43218 10350
rect 43274 10294 43342 10350
rect 43398 10294 60970 10350
rect 61026 10294 61094 10350
rect 61150 10294 61218 10350
rect 61274 10294 61342 10350
rect 61398 10294 78970 10350
rect 79026 10294 79094 10350
rect 79150 10294 79218 10350
rect 79274 10294 79342 10350
rect 79398 10294 96970 10350
rect 97026 10294 97094 10350
rect 97150 10294 97218 10350
rect 97274 10294 97342 10350
rect 97398 10294 114970 10350
rect 115026 10294 115094 10350
rect 115150 10294 115218 10350
rect 115274 10294 115342 10350
rect 115398 10294 132970 10350
rect 133026 10294 133094 10350
rect 133150 10294 133218 10350
rect 133274 10294 133342 10350
rect 133398 10294 150970 10350
rect 151026 10294 151094 10350
rect 151150 10294 151218 10350
rect 151274 10294 151342 10350
rect 151398 10294 168970 10350
rect 169026 10294 169094 10350
rect 169150 10294 169218 10350
rect 169274 10294 169342 10350
rect 169398 10294 186970 10350
rect 187026 10294 187094 10350
rect 187150 10294 187218 10350
rect 187274 10294 187342 10350
rect 187398 10294 204970 10350
rect 205026 10294 205094 10350
rect 205150 10294 205218 10350
rect 205274 10294 205342 10350
rect 205398 10294 222970 10350
rect 223026 10294 223094 10350
rect 223150 10294 223218 10350
rect 223274 10294 223342 10350
rect 223398 10294 240970 10350
rect 241026 10294 241094 10350
rect 241150 10294 241218 10350
rect 241274 10294 241342 10350
rect 241398 10294 258970 10350
rect 259026 10294 259094 10350
rect 259150 10294 259218 10350
rect 259274 10294 259342 10350
rect 259398 10294 276970 10350
rect 277026 10294 277094 10350
rect 277150 10294 277218 10350
rect 277274 10294 277342 10350
rect 277398 10294 294970 10350
rect 295026 10294 295094 10350
rect 295150 10294 295218 10350
rect 295274 10294 295342 10350
rect 295398 10294 312970 10350
rect 313026 10294 313094 10350
rect 313150 10294 313218 10350
rect 313274 10294 313342 10350
rect 313398 10294 330970 10350
rect 331026 10294 331094 10350
rect 331150 10294 331218 10350
rect 331274 10294 331342 10350
rect 331398 10294 348970 10350
rect 349026 10294 349094 10350
rect 349150 10294 349218 10350
rect 349274 10294 349342 10350
rect 349398 10294 366970 10350
rect 367026 10294 367094 10350
rect 367150 10294 367218 10350
rect 367274 10294 367342 10350
rect 367398 10294 384970 10350
rect 385026 10294 385094 10350
rect 385150 10294 385218 10350
rect 385274 10294 385342 10350
rect 385398 10294 402970 10350
rect 403026 10294 403094 10350
rect 403150 10294 403218 10350
rect 403274 10294 403342 10350
rect 403398 10294 420970 10350
rect 421026 10294 421094 10350
rect 421150 10294 421218 10350
rect 421274 10294 421342 10350
rect 421398 10294 438970 10350
rect 439026 10294 439094 10350
rect 439150 10294 439218 10350
rect 439274 10294 439342 10350
rect 439398 10294 456970 10350
rect 457026 10294 457094 10350
rect 457150 10294 457218 10350
rect 457274 10294 457342 10350
rect 457398 10294 474970 10350
rect 475026 10294 475094 10350
rect 475150 10294 475218 10350
rect 475274 10294 475342 10350
rect 475398 10294 492970 10350
rect 493026 10294 493094 10350
rect 493150 10294 493218 10350
rect 493274 10294 493342 10350
rect 493398 10294 510970 10350
rect 511026 10294 511094 10350
rect 511150 10294 511218 10350
rect 511274 10294 511342 10350
rect 511398 10294 528970 10350
rect 529026 10294 529094 10350
rect 529150 10294 529218 10350
rect 529274 10294 529342 10350
rect 529398 10294 546970 10350
rect 547026 10294 547094 10350
rect 547150 10294 547218 10350
rect 547274 10294 547342 10350
rect 547398 10294 564970 10350
rect 565026 10294 565094 10350
rect 565150 10294 565218 10350
rect 565274 10294 565342 10350
rect 565398 10294 582970 10350
rect 583026 10294 583094 10350
rect 583150 10294 583218 10350
rect 583274 10294 583342 10350
rect 583398 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect -1916 10226 597980 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 6970 10226
rect 7026 10170 7094 10226
rect 7150 10170 7218 10226
rect 7274 10170 7342 10226
rect 7398 10170 24970 10226
rect 25026 10170 25094 10226
rect 25150 10170 25218 10226
rect 25274 10170 25342 10226
rect 25398 10170 42970 10226
rect 43026 10170 43094 10226
rect 43150 10170 43218 10226
rect 43274 10170 43342 10226
rect 43398 10170 60970 10226
rect 61026 10170 61094 10226
rect 61150 10170 61218 10226
rect 61274 10170 61342 10226
rect 61398 10170 78970 10226
rect 79026 10170 79094 10226
rect 79150 10170 79218 10226
rect 79274 10170 79342 10226
rect 79398 10170 96970 10226
rect 97026 10170 97094 10226
rect 97150 10170 97218 10226
rect 97274 10170 97342 10226
rect 97398 10170 114970 10226
rect 115026 10170 115094 10226
rect 115150 10170 115218 10226
rect 115274 10170 115342 10226
rect 115398 10170 132970 10226
rect 133026 10170 133094 10226
rect 133150 10170 133218 10226
rect 133274 10170 133342 10226
rect 133398 10170 150970 10226
rect 151026 10170 151094 10226
rect 151150 10170 151218 10226
rect 151274 10170 151342 10226
rect 151398 10170 168970 10226
rect 169026 10170 169094 10226
rect 169150 10170 169218 10226
rect 169274 10170 169342 10226
rect 169398 10170 186970 10226
rect 187026 10170 187094 10226
rect 187150 10170 187218 10226
rect 187274 10170 187342 10226
rect 187398 10170 204970 10226
rect 205026 10170 205094 10226
rect 205150 10170 205218 10226
rect 205274 10170 205342 10226
rect 205398 10170 222970 10226
rect 223026 10170 223094 10226
rect 223150 10170 223218 10226
rect 223274 10170 223342 10226
rect 223398 10170 240970 10226
rect 241026 10170 241094 10226
rect 241150 10170 241218 10226
rect 241274 10170 241342 10226
rect 241398 10170 258970 10226
rect 259026 10170 259094 10226
rect 259150 10170 259218 10226
rect 259274 10170 259342 10226
rect 259398 10170 276970 10226
rect 277026 10170 277094 10226
rect 277150 10170 277218 10226
rect 277274 10170 277342 10226
rect 277398 10170 294970 10226
rect 295026 10170 295094 10226
rect 295150 10170 295218 10226
rect 295274 10170 295342 10226
rect 295398 10170 312970 10226
rect 313026 10170 313094 10226
rect 313150 10170 313218 10226
rect 313274 10170 313342 10226
rect 313398 10170 330970 10226
rect 331026 10170 331094 10226
rect 331150 10170 331218 10226
rect 331274 10170 331342 10226
rect 331398 10170 348970 10226
rect 349026 10170 349094 10226
rect 349150 10170 349218 10226
rect 349274 10170 349342 10226
rect 349398 10170 366970 10226
rect 367026 10170 367094 10226
rect 367150 10170 367218 10226
rect 367274 10170 367342 10226
rect 367398 10170 384970 10226
rect 385026 10170 385094 10226
rect 385150 10170 385218 10226
rect 385274 10170 385342 10226
rect 385398 10170 402970 10226
rect 403026 10170 403094 10226
rect 403150 10170 403218 10226
rect 403274 10170 403342 10226
rect 403398 10170 420970 10226
rect 421026 10170 421094 10226
rect 421150 10170 421218 10226
rect 421274 10170 421342 10226
rect 421398 10170 438970 10226
rect 439026 10170 439094 10226
rect 439150 10170 439218 10226
rect 439274 10170 439342 10226
rect 439398 10170 456970 10226
rect 457026 10170 457094 10226
rect 457150 10170 457218 10226
rect 457274 10170 457342 10226
rect 457398 10170 474970 10226
rect 475026 10170 475094 10226
rect 475150 10170 475218 10226
rect 475274 10170 475342 10226
rect 475398 10170 492970 10226
rect 493026 10170 493094 10226
rect 493150 10170 493218 10226
rect 493274 10170 493342 10226
rect 493398 10170 510970 10226
rect 511026 10170 511094 10226
rect 511150 10170 511218 10226
rect 511274 10170 511342 10226
rect 511398 10170 528970 10226
rect 529026 10170 529094 10226
rect 529150 10170 529218 10226
rect 529274 10170 529342 10226
rect 529398 10170 546970 10226
rect 547026 10170 547094 10226
rect 547150 10170 547218 10226
rect 547274 10170 547342 10226
rect 547398 10170 564970 10226
rect 565026 10170 565094 10226
rect 565150 10170 565218 10226
rect 565274 10170 565342 10226
rect 565398 10170 582970 10226
rect 583026 10170 583094 10226
rect 583150 10170 583218 10226
rect 583274 10170 583342 10226
rect 583398 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect -1916 10102 597980 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 6970 10102
rect 7026 10046 7094 10102
rect 7150 10046 7218 10102
rect 7274 10046 7342 10102
rect 7398 10046 24970 10102
rect 25026 10046 25094 10102
rect 25150 10046 25218 10102
rect 25274 10046 25342 10102
rect 25398 10046 42970 10102
rect 43026 10046 43094 10102
rect 43150 10046 43218 10102
rect 43274 10046 43342 10102
rect 43398 10046 60970 10102
rect 61026 10046 61094 10102
rect 61150 10046 61218 10102
rect 61274 10046 61342 10102
rect 61398 10046 78970 10102
rect 79026 10046 79094 10102
rect 79150 10046 79218 10102
rect 79274 10046 79342 10102
rect 79398 10046 96970 10102
rect 97026 10046 97094 10102
rect 97150 10046 97218 10102
rect 97274 10046 97342 10102
rect 97398 10046 114970 10102
rect 115026 10046 115094 10102
rect 115150 10046 115218 10102
rect 115274 10046 115342 10102
rect 115398 10046 132970 10102
rect 133026 10046 133094 10102
rect 133150 10046 133218 10102
rect 133274 10046 133342 10102
rect 133398 10046 150970 10102
rect 151026 10046 151094 10102
rect 151150 10046 151218 10102
rect 151274 10046 151342 10102
rect 151398 10046 168970 10102
rect 169026 10046 169094 10102
rect 169150 10046 169218 10102
rect 169274 10046 169342 10102
rect 169398 10046 186970 10102
rect 187026 10046 187094 10102
rect 187150 10046 187218 10102
rect 187274 10046 187342 10102
rect 187398 10046 204970 10102
rect 205026 10046 205094 10102
rect 205150 10046 205218 10102
rect 205274 10046 205342 10102
rect 205398 10046 222970 10102
rect 223026 10046 223094 10102
rect 223150 10046 223218 10102
rect 223274 10046 223342 10102
rect 223398 10046 240970 10102
rect 241026 10046 241094 10102
rect 241150 10046 241218 10102
rect 241274 10046 241342 10102
rect 241398 10046 258970 10102
rect 259026 10046 259094 10102
rect 259150 10046 259218 10102
rect 259274 10046 259342 10102
rect 259398 10046 276970 10102
rect 277026 10046 277094 10102
rect 277150 10046 277218 10102
rect 277274 10046 277342 10102
rect 277398 10046 294970 10102
rect 295026 10046 295094 10102
rect 295150 10046 295218 10102
rect 295274 10046 295342 10102
rect 295398 10046 312970 10102
rect 313026 10046 313094 10102
rect 313150 10046 313218 10102
rect 313274 10046 313342 10102
rect 313398 10046 330970 10102
rect 331026 10046 331094 10102
rect 331150 10046 331218 10102
rect 331274 10046 331342 10102
rect 331398 10046 348970 10102
rect 349026 10046 349094 10102
rect 349150 10046 349218 10102
rect 349274 10046 349342 10102
rect 349398 10046 366970 10102
rect 367026 10046 367094 10102
rect 367150 10046 367218 10102
rect 367274 10046 367342 10102
rect 367398 10046 384970 10102
rect 385026 10046 385094 10102
rect 385150 10046 385218 10102
rect 385274 10046 385342 10102
rect 385398 10046 402970 10102
rect 403026 10046 403094 10102
rect 403150 10046 403218 10102
rect 403274 10046 403342 10102
rect 403398 10046 420970 10102
rect 421026 10046 421094 10102
rect 421150 10046 421218 10102
rect 421274 10046 421342 10102
rect 421398 10046 438970 10102
rect 439026 10046 439094 10102
rect 439150 10046 439218 10102
rect 439274 10046 439342 10102
rect 439398 10046 456970 10102
rect 457026 10046 457094 10102
rect 457150 10046 457218 10102
rect 457274 10046 457342 10102
rect 457398 10046 474970 10102
rect 475026 10046 475094 10102
rect 475150 10046 475218 10102
rect 475274 10046 475342 10102
rect 475398 10046 492970 10102
rect 493026 10046 493094 10102
rect 493150 10046 493218 10102
rect 493274 10046 493342 10102
rect 493398 10046 510970 10102
rect 511026 10046 511094 10102
rect 511150 10046 511218 10102
rect 511274 10046 511342 10102
rect 511398 10046 528970 10102
rect 529026 10046 529094 10102
rect 529150 10046 529218 10102
rect 529274 10046 529342 10102
rect 529398 10046 546970 10102
rect 547026 10046 547094 10102
rect 547150 10046 547218 10102
rect 547274 10046 547342 10102
rect 547398 10046 564970 10102
rect 565026 10046 565094 10102
rect 565150 10046 565218 10102
rect 565274 10046 565342 10102
rect 565398 10046 582970 10102
rect 583026 10046 583094 10102
rect 583150 10046 583218 10102
rect 583274 10046 583342 10102
rect 583398 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect -1916 9978 597980 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 6970 9978
rect 7026 9922 7094 9978
rect 7150 9922 7218 9978
rect 7274 9922 7342 9978
rect 7398 9922 24970 9978
rect 25026 9922 25094 9978
rect 25150 9922 25218 9978
rect 25274 9922 25342 9978
rect 25398 9922 42970 9978
rect 43026 9922 43094 9978
rect 43150 9922 43218 9978
rect 43274 9922 43342 9978
rect 43398 9922 60970 9978
rect 61026 9922 61094 9978
rect 61150 9922 61218 9978
rect 61274 9922 61342 9978
rect 61398 9922 78970 9978
rect 79026 9922 79094 9978
rect 79150 9922 79218 9978
rect 79274 9922 79342 9978
rect 79398 9922 96970 9978
rect 97026 9922 97094 9978
rect 97150 9922 97218 9978
rect 97274 9922 97342 9978
rect 97398 9922 114970 9978
rect 115026 9922 115094 9978
rect 115150 9922 115218 9978
rect 115274 9922 115342 9978
rect 115398 9922 132970 9978
rect 133026 9922 133094 9978
rect 133150 9922 133218 9978
rect 133274 9922 133342 9978
rect 133398 9922 150970 9978
rect 151026 9922 151094 9978
rect 151150 9922 151218 9978
rect 151274 9922 151342 9978
rect 151398 9922 168970 9978
rect 169026 9922 169094 9978
rect 169150 9922 169218 9978
rect 169274 9922 169342 9978
rect 169398 9922 186970 9978
rect 187026 9922 187094 9978
rect 187150 9922 187218 9978
rect 187274 9922 187342 9978
rect 187398 9922 204970 9978
rect 205026 9922 205094 9978
rect 205150 9922 205218 9978
rect 205274 9922 205342 9978
rect 205398 9922 222970 9978
rect 223026 9922 223094 9978
rect 223150 9922 223218 9978
rect 223274 9922 223342 9978
rect 223398 9922 240970 9978
rect 241026 9922 241094 9978
rect 241150 9922 241218 9978
rect 241274 9922 241342 9978
rect 241398 9922 258970 9978
rect 259026 9922 259094 9978
rect 259150 9922 259218 9978
rect 259274 9922 259342 9978
rect 259398 9922 276970 9978
rect 277026 9922 277094 9978
rect 277150 9922 277218 9978
rect 277274 9922 277342 9978
rect 277398 9922 294970 9978
rect 295026 9922 295094 9978
rect 295150 9922 295218 9978
rect 295274 9922 295342 9978
rect 295398 9922 312970 9978
rect 313026 9922 313094 9978
rect 313150 9922 313218 9978
rect 313274 9922 313342 9978
rect 313398 9922 330970 9978
rect 331026 9922 331094 9978
rect 331150 9922 331218 9978
rect 331274 9922 331342 9978
rect 331398 9922 348970 9978
rect 349026 9922 349094 9978
rect 349150 9922 349218 9978
rect 349274 9922 349342 9978
rect 349398 9922 366970 9978
rect 367026 9922 367094 9978
rect 367150 9922 367218 9978
rect 367274 9922 367342 9978
rect 367398 9922 384970 9978
rect 385026 9922 385094 9978
rect 385150 9922 385218 9978
rect 385274 9922 385342 9978
rect 385398 9922 402970 9978
rect 403026 9922 403094 9978
rect 403150 9922 403218 9978
rect 403274 9922 403342 9978
rect 403398 9922 420970 9978
rect 421026 9922 421094 9978
rect 421150 9922 421218 9978
rect 421274 9922 421342 9978
rect 421398 9922 438970 9978
rect 439026 9922 439094 9978
rect 439150 9922 439218 9978
rect 439274 9922 439342 9978
rect 439398 9922 456970 9978
rect 457026 9922 457094 9978
rect 457150 9922 457218 9978
rect 457274 9922 457342 9978
rect 457398 9922 474970 9978
rect 475026 9922 475094 9978
rect 475150 9922 475218 9978
rect 475274 9922 475342 9978
rect 475398 9922 492970 9978
rect 493026 9922 493094 9978
rect 493150 9922 493218 9978
rect 493274 9922 493342 9978
rect 493398 9922 510970 9978
rect 511026 9922 511094 9978
rect 511150 9922 511218 9978
rect 511274 9922 511342 9978
rect 511398 9922 528970 9978
rect 529026 9922 529094 9978
rect 529150 9922 529218 9978
rect 529274 9922 529342 9978
rect 529398 9922 546970 9978
rect 547026 9922 547094 9978
rect 547150 9922 547218 9978
rect 547274 9922 547342 9978
rect 547398 9922 564970 9978
rect 565026 9922 565094 9978
rect 565150 9922 565218 9978
rect 565274 9922 565342 9978
rect 565398 9922 582970 9978
rect 583026 9922 583094 9978
rect 583150 9922 583218 9978
rect 583274 9922 583342 9978
rect 583398 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect -1916 9826 597980 9922
rect -1916 4350 597980 4446
rect -1916 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 3250 4350
rect 3306 4294 3374 4350
rect 3430 4294 3498 4350
rect 3554 4294 3622 4350
rect 3678 4294 21250 4350
rect 21306 4294 21374 4350
rect 21430 4294 21498 4350
rect 21554 4294 21622 4350
rect 21678 4294 39250 4350
rect 39306 4294 39374 4350
rect 39430 4294 39498 4350
rect 39554 4294 39622 4350
rect 39678 4294 57250 4350
rect 57306 4294 57374 4350
rect 57430 4294 57498 4350
rect 57554 4294 57622 4350
rect 57678 4294 75250 4350
rect 75306 4294 75374 4350
rect 75430 4294 75498 4350
rect 75554 4294 75622 4350
rect 75678 4294 93250 4350
rect 93306 4294 93374 4350
rect 93430 4294 93498 4350
rect 93554 4294 93622 4350
rect 93678 4294 111250 4350
rect 111306 4294 111374 4350
rect 111430 4294 111498 4350
rect 111554 4294 111622 4350
rect 111678 4294 129250 4350
rect 129306 4294 129374 4350
rect 129430 4294 129498 4350
rect 129554 4294 129622 4350
rect 129678 4294 147250 4350
rect 147306 4294 147374 4350
rect 147430 4294 147498 4350
rect 147554 4294 147622 4350
rect 147678 4294 165250 4350
rect 165306 4294 165374 4350
rect 165430 4294 165498 4350
rect 165554 4294 165622 4350
rect 165678 4294 183250 4350
rect 183306 4294 183374 4350
rect 183430 4294 183498 4350
rect 183554 4294 183622 4350
rect 183678 4294 201250 4350
rect 201306 4294 201374 4350
rect 201430 4294 201498 4350
rect 201554 4294 201622 4350
rect 201678 4294 219250 4350
rect 219306 4294 219374 4350
rect 219430 4294 219498 4350
rect 219554 4294 219622 4350
rect 219678 4294 237250 4350
rect 237306 4294 237374 4350
rect 237430 4294 237498 4350
rect 237554 4294 237622 4350
rect 237678 4294 255250 4350
rect 255306 4294 255374 4350
rect 255430 4294 255498 4350
rect 255554 4294 255622 4350
rect 255678 4294 273250 4350
rect 273306 4294 273374 4350
rect 273430 4294 273498 4350
rect 273554 4294 273622 4350
rect 273678 4294 291250 4350
rect 291306 4294 291374 4350
rect 291430 4294 291498 4350
rect 291554 4294 291622 4350
rect 291678 4294 309250 4350
rect 309306 4294 309374 4350
rect 309430 4294 309498 4350
rect 309554 4294 309622 4350
rect 309678 4294 327250 4350
rect 327306 4294 327374 4350
rect 327430 4294 327498 4350
rect 327554 4294 327622 4350
rect 327678 4294 345250 4350
rect 345306 4294 345374 4350
rect 345430 4294 345498 4350
rect 345554 4294 345622 4350
rect 345678 4294 363250 4350
rect 363306 4294 363374 4350
rect 363430 4294 363498 4350
rect 363554 4294 363622 4350
rect 363678 4294 381250 4350
rect 381306 4294 381374 4350
rect 381430 4294 381498 4350
rect 381554 4294 381622 4350
rect 381678 4294 399250 4350
rect 399306 4294 399374 4350
rect 399430 4294 399498 4350
rect 399554 4294 399622 4350
rect 399678 4294 417250 4350
rect 417306 4294 417374 4350
rect 417430 4294 417498 4350
rect 417554 4294 417622 4350
rect 417678 4294 435250 4350
rect 435306 4294 435374 4350
rect 435430 4294 435498 4350
rect 435554 4294 435622 4350
rect 435678 4294 453250 4350
rect 453306 4294 453374 4350
rect 453430 4294 453498 4350
rect 453554 4294 453622 4350
rect 453678 4294 471250 4350
rect 471306 4294 471374 4350
rect 471430 4294 471498 4350
rect 471554 4294 471622 4350
rect 471678 4294 489250 4350
rect 489306 4294 489374 4350
rect 489430 4294 489498 4350
rect 489554 4294 489622 4350
rect 489678 4294 507250 4350
rect 507306 4294 507374 4350
rect 507430 4294 507498 4350
rect 507554 4294 507622 4350
rect 507678 4294 525250 4350
rect 525306 4294 525374 4350
rect 525430 4294 525498 4350
rect 525554 4294 525622 4350
rect 525678 4294 543250 4350
rect 543306 4294 543374 4350
rect 543430 4294 543498 4350
rect 543554 4294 543622 4350
rect 543678 4294 561250 4350
rect 561306 4294 561374 4350
rect 561430 4294 561498 4350
rect 561554 4294 561622 4350
rect 561678 4294 579250 4350
rect 579306 4294 579374 4350
rect 579430 4294 579498 4350
rect 579554 4294 579622 4350
rect 579678 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597980 4350
rect -1916 4226 597980 4294
rect -1916 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 3250 4226
rect 3306 4170 3374 4226
rect 3430 4170 3498 4226
rect 3554 4170 3622 4226
rect 3678 4170 21250 4226
rect 21306 4170 21374 4226
rect 21430 4170 21498 4226
rect 21554 4170 21622 4226
rect 21678 4170 39250 4226
rect 39306 4170 39374 4226
rect 39430 4170 39498 4226
rect 39554 4170 39622 4226
rect 39678 4170 57250 4226
rect 57306 4170 57374 4226
rect 57430 4170 57498 4226
rect 57554 4170 57622 4226
rect 57678 4170 75250 4226
rect 75306 4170 75374 4226
rect 75430 4170 75498 4226
rect 75554 4170 75622 4226
rect 75678 4170 93250 4226
rect 93306 4170 93374 4226
rect 93430 4170 93498 4226
rect 93554 4170 93622 4226
rect 93678 4170 111250 4226
rect 111306 4170 111374 4226
rect 111430 4170 111498 4226
rect 111554 4170 111622 4226
rect 111678 4170 129250 4226
rect 129306 4170 129374 4226
rect 129430 4170 129498 4226
rect 129554 4170 129622 4226
rect 129678 4170 147250 4226
rect 147306 4170 147374 4226
rect 147430 4170 147498 4226
rect 147554 4170 147622 4226
rect 147678 4170 165250 4226
rect 165306 4170 165374 4226
rect 165430 4170 165498 4226
rect 165554 4170 165622 4226
rect 165678 4170 183250 4226
rect 183306 4170 183374 4226
rect 183430 4170 183498 4226
rect 183554 4170 183622 4226
rect 183678 4170 201250 4226
rect 201306 4170 201374 4226
rect 201430 4170 201498 4226
rect 201554 4170 201622 4226
rect 201678 4170 219250 4226
rect 219306 4170 219374 4226
rect 219430 4170 219498 4226
rect 219554 4170 219622 4226
rect 219678 4170 237250 4226
rect 237306 4170 237374 4226
rect 237430 4170 237498 4226
rect 237554 4170 237622 4226
rect 237678 4170 255250 4226
rect 255306 4170 255374 4226
rect 255430 4170 255498 4226
rect 255554 4170 255622 4226
rect 255678 4170 273250 4226
rect 273306 4170 273374 4226
rect 273430 4170 273498 4226
rect 273554 4170 273622 4226
rect 273678 4170 291250 4226
rect 291306 4170 291374 4226
rect 291430 4170 291498 4226
rect 291554 4170 291622 4226
rect 291678 4170 309250 4226
rect 309306 4170 309374 4226
rect 309430 4170 309498 4226
rect 309554 4170 309622 4226
rect 309678 4170 327250 4226
rect 327306 4170 327374 4226
rect 327430 4170 327498 4226
rect 327554 4170 327622 4226
rect 327678 4170 345250 4226
rect 345306 4170 345374 4226
rect 345430 4170 345498 4226
rect 345554 4170 345622 4226
rect 345678 4170 363250 4226
rect 363306 4170 363374 4226
rect 363430 4170 363498 4226
rect 363554 4170 363622 4226
rect 363678 4170 381250 4226
rect 381306 4170 381374 4226
rect 381430 4170 381498 4226
rect 381554 4170 381622 4226
rect 381678 4170 399250 4226
rect 399306 4170 399374 4226
rect 399430 4170 399498 4226
rect 399554 4170 399622 4226
rect 399678 4170 417250 4226
rect 417306 4170 417374 4226
rect 417430 4170 417498 4226
rect 417554 4170 417622 4226
rect 417678 4170 435250 4226
rect 435306 4170 435374 4226
rect 435430 4170 435498 4226
rect 435554 4170 435622 4226
rect 435678 4170 453250 4226
rect 453306 4170 453374 4226
rect 453430 4170 453498 4226
rect 453554 4170 453622 4226
rect 453678 4170 471250 4226
rect 471306 4170 471374 4226
rect 471430 4170 471498 4226
rect 471554 4170 471622 4226
rect 471678 4170 489250 4226
rect 489306 4170 489374 4226
rect 489430 4170 489498 4226
rect 489554 4170 489622 4226
rect 489678 4170 507250 4226
rect 507306 4170 507374 4226
rect 507430 4170 507498 4226
rect 507554 4170 507622 4226
rect 507678 4170 525250 4226
rect 525306 4170 525374 4226
rect 525430 4170 525498 4226
rect 525554 4170 525622 4226
rect 525678 4170 543250 4226
rect 543306 4170 543374 4226
rect 543430 4170 543498 4226
rect 543554 4170 543622 4226
rect 543678 4170 561250 4226
rect 561306 4170 561374 4226
rect 561430 4170 561498 4226
rect 561554 4170 561622 4226
rect 561678 4170 579250 4226
rect 579306 4170 579374 4226
rect 579430 4170 579498 4226
rect 579554 4170 579622 4226
rect 579678 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597980 4226
rect -1916 4102 597980 4170
rect -1916 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 3250 4102
rect 3306 4046 3374 4102
rect 3430 4046 3498 4102
rect 3554 4046 3622 4102
rect 3678 4046 21250 4102
rect 21306 4046 21374 4102
rect 21430 4046 21498 4102
rect 21554 4046 21622 4102
rect 21678 4046 39250 4102
rect 39306 4046 39374 4102
rect 39430 4046 39498 4102
rect 39554 4046 39622 4102
rect 39678 4046 57250 4102
rect 57306 4046 57374 4102
rect 57430 4046 57498 4102
rect 57554 4046 57622 4102
rect 57678 4046 75250 4102
rect 75306 4046 75374 4102
rect 75430 4046 75498 4102
rect 75554 4046 75622 4102
rect 75678 4046 93250 4102
rect 93306 4046 93374 4102
rect 93430 4046 93498 4102
rect 93554 4046 93622 4102
rect 93678 4046 111250 4102
rect 111306 4046 111374 4102
rect 111430 4046 111498 4102
rect 111554 4046 111622 4102
rect 111678 4046 129250 4102
rect 129306 4046 129374 4102
rect 129430 4046 129498 4102
rect 129554 4046 129622 4102
rect 129678 4046 147250 4102
rect 147306 4046 147374 4102
rect 147430 4046 147498 4102
rect 147554 4046 147622 4102
rect 147678 4046 165250 4102
rect 165306 4046 165374 4102
rect 165430 4046 165498 4102
rect 165554 4046 165622 4102
rect 165678 4046 183250 4102
rect 183306 4046 183374 4102
rect 183430 4046 183498 4102
rect 183554 4046 183622 4102
rect 183678 4046 201250 4102
rect 201306 4046 201374 4102
rect 201430 4046 201498 4102
rect 201554 4046 201622 4102
rect 201678 4046 219250 4102
rect 219306 4046 219374 4102
rect 219430 4046 219498 4102
rect 219554 4046 219622 4102
rect 219678 4046 237250 4102
rect 237306 4046 237374 4102
rect 237430 4046 237498 4102
rect 237554 4046 237622 4102
rect 237678 4046 255250 4102
rect 255306 4046 255374 4102
rect 255430 4046 255498 4102
rect 255554 4046 255622 4102
rect 255678 4046 273250 4102
rect 273306 4046 273374 4102
rect 273430 4046 273498 4102
rect 273554 4046 273622 4102
rect 273678 4046 291250 4102
rect 291306 4046 291374 4102
rect 291430 4046 291498 4102
rect 291554 4046 291622 4102
rect 291678 4046 309250 4102
rect 309306 4046 309374 4102
rect 309430 4046 309498 4102
rect 309554 4046 309622 4102
rect 309678 4046 327250 4102
rect 327306 4046 327374 4102
rect 327430 4046 327498 4102
rect 327554 4046 327622 4102
rect 327678 4046 345250 4102
rect 345306 4046 345374 4102
rect 345430 4046 345498 4102
rect 345554 4046 345622 4102
rect 345678 4046 363250 4102
rect 363306 4046 363374 4102
rect 363430 4046 363498 4102
rect 363554 4046 363622 4102
rect 363678 4046 381250 4102
rect 381306 4046 381374 4102
rect 381430 4046 381498 4102
rect 381554 4046 381622 4102
rect 381678 4046 399250 4102
rect 399306 4046 399374 4102
rect 399430 4046 399498 4102
rect 399554 4046 399622 4102
rect 399678 4046 417250 4102
rect 417306 4046 417374 4102
rect 417430 4046 417498 4102
rect 417554 4046 417622 4102
rect 417678 4046 435250 4102
rect 435306 4046 435374 4102
rect 435430 4046 435498 4102
rect 435554 4046 435622 4102
rect 435678 4046 453250 4102
rect 453306 4046 453374 4102
rect 453430 4046 453498 4102
rect 453554 4046 453622 4102
rect 453678 4046 471250 4102
rect 471306 4046 471374 4102
rect 471430 4046 471498 4102
rect 471554 4046 471622 4102
rect 471678 4046 489250 4102
rect 489306 4046 489374 4102
rect 489430 4046 489498 4102
rect 489554 4046 489622 4102
rect 489678 4046 507250 4102
rect 507306 4046 507374 4102
rect 507430 4046 507498 4102
rect 507554 4046 507622 4102
rect 507678 4046 525250 4102
rect 525306 4046 525374 4102
rect 525430 4046 525498 4102
rect 525554 4046 525622 4102
rect 525678 4046 543250 4102
rect 543306 4046 543374 4102
rect 543430 4046 543498 4102
rect 543554 4046 543622 4102
rect 543678 4046 561250 4102
rect 561306 4046 561374 4102
rect 561430 4046 561498 4102
rect 561554 4046 561622 4102
rect 561678 4046 579250 4102
rect 579306 4046 579374 4102
rect 579430 4046 579498 4102
rect 579554 4046 579622 4102
rect 579678 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597980 4102
rect -1916 3978 597980 4046
rect -1916 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 3250 3978
rect 3306 3922 3374 3978
rect 3430 3922 3498 3978
rect 3554 3922 3622 3978
rect 3678 3922 21250 3978
rect 21306 3922 21374 3978
rect 21430 3922 21498 3978
rect 21554 3922 21622 3978
rect 21678 3922 39250 3978
rect 39306 3922 39374 3978
rect 39430 3922 39498 3978
rect 39554 3922 39622 3978
rect 39678 3922 57250 3978
rect 57306 3922 57374 3978
rect 57430 3922 57498 3978
rect 57554 3922 57622 3978
rect 57678 3922 75250 3978
rect 75306 3922 75374 3978
rect 75430 3922 75498 3978
rect 75554 3922 75622 3978
rect 75678 3922 93250 3978
rect 93306 3922 93374 3978
rect 93430 3922 93498 3978
rect 93554 3922 93622 3978
rect 93678 3922 111250 3978
rect 111306 3922 111374 3978
rect 111430 3922 111498 3978
rect 111554 3922 111622 3978
rect 111678 3922 129250 3978
rect 129306 3922 129374 3978
rect 129430 3922 129498 3978
rect 129554 3922 129622 3978
rect 129678 3922 147250 3978
rect 147306 3922 147374 3978
rect 147430 3922 147498 3978
rect 147554 3922 147622 3978
rect 147678 3922 165250 3978
rect 165306 3922 165374 3978
rect 165430 3922 165498 3978
rect 165554 3922 165622 3978
rect 165678 3922 183250 3978
rect 183306 3922 183374 3978
rect 183430 3922 183498 3978
rect 183554 3922 183622 3978
rect 183678 3922 201250 3978
rect 201306 3922 201374 3978
rect 201430 3922 201498 3978
rect 201554 3922 201622 3978
rect 201678 3922 219250 3978
rect 219306 3922 219374 3978
rect 219430 3922 219498 3978
rect 219554 3922 219622 3978
rect 219678 3922 237250 3978
rect 237306 3922 237374 3978
rect 237430 3922 237498 3978
rect 237554 3922 237622 3978
rect 237678 3922 255250 3978
rect 255306 3922 255374 3978
rect 255430 3922 255498 3978
rect 255554 3922 255622 3978
rect 255678 3922 273250 3978
rect 273306 3922 273374 3978
rect 273430 3922 273498 3978
rect 273554 3922 273622 3978
rect 273678 3922 291250 3978
rect 291306 3922 291374 3978
rect 291430 3922 291498 3978
rect 291554 3922 291622 3978
rect 291678 3922 309250 3978
rect 309306 3922 309374 3978
rect 309430 3922 309498 3978
rect 309554 3922 309622 3978
rect 309678 3922 327250 3978
rect 327306 3922 327374 3978
rect 327430 3922 327498 3978
rect 327554 3922 327622 3978
rect 327678 3922 345250 3978
rect 345306 3922 345374 3978
rect 345430 3922 345498 3978
rect 345554 3922 345622 3978
rect 345678 3922 363250 3978
rect 363306 3922 363374 3978
rect 363430 3922 363498 3978
rect 363554 3922 363622 3978
rect 363678 3922 381250 3978
rect 381306 3922 381374 3978
rect 381430 3922 381498 3978
rect 381554 3922 381622 3978
rect 381678 3922 399250 3978
rect 399306 3922 399374 3978
rect 399430 3922 399498 3978
rect 399554 3922 399622 3978
rect 399678 3922 417250 3978
rect 417306 3922 417374 3978
rect 417430 3922 417498 3978
rect 417554 3922 417622 3978
rect 417678 3922 435250 3978
rect 435306 3922 435374 3978
rect 435430 3922 435498 3978
rect 435554 3922 435622 3978
rect 435678 3922 453250 3978
rect 453306 3922 453374 3978
rect 453430 3922 453498 3978
rect 453554 3922 453622 3978
rect 453678 3922 471250 3978
rect 471306 3922 471374 3978
rect 471430 3922 471498 3978
rect 471554 3922 471622 3978
rect 471678 3922 489250 3978
rect 489306 3922 489374 3978
rect 489430 3922 489498 3978
rect 489554 3922 489622 3978
rect 489678 3922 507250 3978
rect 507306 3922 507374 3978
rect 507430 3922 507498 3978
rect 507554 3922 507622 3978
rect 507678 3922 525250 3978
rect 525306 3922 525374 3978
rect 525430 3922 525498 3978
rect 525554 3922 525622 3978
rect 525678 3922 543250 3978
rect 543306 3922 543374 3978
rect 543430 3922 543498 3978
rect 543554 3922 543622 3978
rect 543678 3922 561250 3978
rect 561306 3922 561374 3978
rect 561430 3922 561498 3978
rect 561554 3922 561622 3978
rect 561678 3922 579250 3978
rect 579306 3922 579374 3978
rect 579430 3922 579498 3978
rect 579554 3922 579622 3978
rect 579678 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597980 3978
rect -1916 3826 597980 3922
rect -956 -160 597020 -64
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 3250 -160
rect 3306 -216 3374 -160
rect 3430 -216 3498 -160
rect 3554 -216 3622 -160
rect 3678 -216 21250 -160
rect 21306 -216 21374 -160
rect 21430 -216 21498 -160
rect 21554 -216 21622 -160
rect 21678 -216 39250 -160
rect 39306 -216 39374 -160
rect 39430 -216 39498 -160
rect 39554 -216 39622 -160
rect 39678 -216 57250 -160
rect 57306 -216 57374 -160
rect 57430 -216 57498 -160
rect 57554 -216 57622 -160
rect 57678 -216 75250 -160
rect 75306 -216 75374 -160
rect 75430 -216 75498 -160
rect 75554 -216 75622 -160
rect 75678 -216 93250 -160
rect 93306 -216 93374 -160
rect 93430 -216 93498 -160
rect 93554 -216 93622 -160
rect 93678 -216 111250 -160
rect 111306 -216 111374 -160
rect 111430 -216 111498 -160
rect 111554 -216 111622 -160
rect 111678 -216 129250 -160
rect 129306 -216 129374 -160
rect 129430 -216 129498 -160
rect 129554 -216 129622 -160
rect 129678 -216 147250 -160
rect 147306 -216 147374 -160
rect 147430 -216 147498 -160
rect 147554 -216 147622 -160
rect 147678 -216 165250 -160
rect 165306 -216 165374 -160
rect 165430 -216 165498 -160
rect 165554 -216 165622 -160
rect 165678 -216 183250 -160
rect 183306 -216 183374 -160
rect 183430 -216 183498 -160
rect 183554 -216 183622 -160
rect 183678 -216 201250 -160
rect 201306 -216 201374 -160
rect 201430 -216 201498 -160
rect 201554 -216 201622 -160
rect 201678 -216 219250 -160
rect 219306 -216 219374 -160
rect 219430 -216 219498 -160
rect 219554 -216 219622 -160
rect 219678 -216 237250 -160
rect 237306 -216 237374 -160
rect 237430 -216 237498 -160
rect 237554 -216 237622 -160
rect 237678 -216 255250 -160
rect 255306 -216 255374 -160
rect 255430 -216 255498 -160
rect 255554 -216 255622 -160
rect 255678 -216 273250 -160
rect 273306 -216 273374 -160
rect 273430 -216 273498 -160
rect 273554 -216 273622 -160
rect 273678 -216 291250 -160
rect 291306 -216 291374 -160
rect 291430 -216 291498 -160
rect 291554 -216 291622 -160
rect 291678 -216 309250 -160
rect 309306 -216 309374 -160
rect 309430 -216 309498 -160
rect 309554 -216 309622 -160
rect 309678 -216 327250 -160
rect 327306 -216 327374 -160
rect 327430 -216 327498 -160
rect 327554 -216 327622 -160
rect 327678 -216 345250 -160
rect 345306 -216 345374 -160
rect 345430 -216 345498 -160
rect 345554 -216 345622 -160
rect 345678 -216 363250 -160
rect 363306 -216 363374 -160
rect 363430 -216 363498 -160
rect 363554 -216 363622 -160
rect 363678 -216 381250 -160
rect 381306 -216 381374 -160
rect 381430 -216 381498 -160
rect 381554 -216 381622 -160
rect 381678 -216 399250 -160
rect 399306 -216 399374 -160
rect 399430 -216 399498 -160
rect 399554 -216 399622 -160
rect 399678 -216 417250 -160
rect 417306 -216 417374 -160
rect 417430 -216 417498 -160
rect 417554 -216 417622 -160
rect 417678 -216 435250 -160
rect 435306 -216 435374 -160
rect 435430 -216 435498 -160
rect 435554 -216 435622 -160
rect 435678 -216 453250 -160
rect 453306 -216 453374 -160
rect 453430 -216 453498 -160
rect 453554 -216 453622 -160
rect 453678 -216 471250 -160
rect 471306 -216 471374 -160
rect 471430 -216 471498 -160
rect 471554 -216 471622 -160
rect 471678 -216 489250 -160
rect 489306 -216 489374 -160
rect 489430 -216 489498 -160
rect 489554 -216 489622 -160
rect 489678 -216 507250 -160
rect 507306 -216 507374 -160
rect 507430 -216 507498 -160
rect 507554 -216 507622 -160
rect 507678 -216 525250 -160
rect 525306 -216 525374 -160
rect 525430 -216 525498 -160
rect 525554 -216 525622 -160
rect 525678 -216 543250 -160
rect 543306 -216 543374 -160
rect 543430 -216 543498 -160
rect 543554 -216 543622 -160
rect 543678 -216 561250 -160
rect 561306 -216 561374 -160
rect 561430 -216 561498 -160
rect 561554 -216 561622 -160
rect 561678 -216 579250 -160
rect 579306 -216 579374 -160
rect 579430 -216 579498 -160
rect 579554 -216 579622 -160
rect 579678 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect -956 -284 597020 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 3250 -284
rect 3306 -340 3374 -284
rect 3430 -340 3498 -284
rect 3554 -340 3622 -284
rect 3678 -340 21250 -284
rect 21306 -340 21374 -284
rect 21430 -340 21498 -284
rect 21554 -340 21622 -284
rect 21678 -340 39250 -284
rect 39306 -340 39374 -284
rect 39430 -340 39498 -284
rect 39554 -340 39622 -284
rect 39678 -340 57250 -284
rect 57306 -340 57374 -284
rect 57430 -340 57498 -284
rect 57554 -340 57622 -284
rect 57678 -340 75250 -284
rect 75306 -340 75374 -284
rect 75430 -340 75498 -284
rect 75554 -340 75622 -284
rect 75678 -340 93250 -284
rect 93306 -340 93374 -284
rect 93430 -340 93498 -284
rect 93554 -340 93622 -284
rect 93678 -340 111250 -284
rect 111306 -340 111374 -284
rect 111430 -340 111498 -284
rect 111554 -340 111622 -284
rect 111678 -340 129250 -284
rect 129306 -340 129374 -284
rect 129430 -340 129498 -284
rect 129554 -340 129622 -284
rect 129678 -340 147250 -284
rect 147306 -340 147374 -284
rect 147430 -340 147498 -284
rect 147554 -340 147622 -284
rect 147678 -340 165250 -284
rect 165306 -340 165374 -284
rect 165430 -340 165498 -284
rect 165554 -340 165622 -284
rect 165678 -340 183250 -284
rect 183306 -340 183374 -284
rect 183430 -340 183498 -284
rect 183554 -340 183622 -284
rect 183678 -340 201250 -284
rect 201306 -340 201374 -284
rect 201430 -340 201498 -284
rect 201554 -340 201622 -284
rect 201678 -340 219250 -284
rect 219306 -340 219374 -284
rect 219430 -340 219498 -284
rect 219554 -340 219622 -284
rect 219678 -340 237250 -284
rect 237306 -340 237374 -284
rect 237430 -340 237498 -284
rect 237554 -340 237622 -284
rect 237678 -340 255250 -284
rect 255306 -340 255374 -284
rect 255430 -340 255498 -284
rect 255554 -340 255622 -284
rect 255678 -340 273250 -284
rect 273306 -340 273374 -284
rect 273430 -340 273498 -284
rect 273554 -340 273622 -284
rect 273678 -340 291250 -284
rect 291306 -340 291374 -284
rect 291430 -340 291498 -284
rect 291554 -340 291622 -284
rect 291678 -340 309250 -284
rect 309306 -340 309374 -284
rect 309430 -340 309498 -284
rect 309554 -340 309622 -284
rect 309678 -340 327250 -284
rect 327306 -340 327374 -284
rect 327430 -340 327498 -284
rect 327554 -340 327622 -284
rect 327678 -340 345250 -284
rect 345306 -340 345374 -284
rect 345430 -340 345498 -284
rect 345554 -340 345622 -284
rect 345678 -340 363250 -284
rect 363306 -340 363374 -284
rect 363430 -340 363498 -284
rect 363554 -340 363622 -284
rect 363678 -340 381250 -284
rect 381306 -340 381374 -284
rect 381430 -340 381498 -284
rect 381554 -340 381622 -284
rect 381678 -340 399250 -284
rect 399306 -340 399374 -284
rect 399430 -340 399498 -284
rect 399554 -340 399622 -284
rect 399678 -340 417250 -284
rect 417306 -340 417374 -284
rect 417430 -340 417498 -284
rect 417554 -340 417622 -284
rect 417678 -340 435250 -284
rect 435306 -340 435374 -284
rect 435430 -340 435498 -284
rect 435554 -340 435622 -284
rect 435678 -340 453250 -284
rect 453306 -340 453374 -284
rect 453430 -340 453498 -284
rect 453554 -340 453622 -284
rect 453678 -340 471250 -284
rect 471306 -340 471374 -284
rect 471430 -340 471498 -284
rect 471554 -340 471622 -284
rect 471678 -340 489250 -284
rect 489306 -340 489374 -284
rect 489430 -340 489498 -284
rect 489554 -340 489622 -284
rect 489678 -340 507250 -284
rect 507306 -340 507374 -284
rect 507430 -340 507498 -284
rect 507554 -340 507622 -284
rect 507678 -340 525250 -284
rect 525306 -340 525374 -284
rect 525430 -340 525498 -284
rect 525554 -340 525622 -284
rect 525678 -340 543250 -284
rect 543306 -340 543374 -284
rect 543430 -340 543498 -284
rect 543554 -340 543622 -284
rect 543678 -340 561250 -284
rect 561306 -340 561374 -284
rect 561430 -340 561498 -284
rect 561554 -340 561622 -284
rect 561678 -340 579250 -284
rect 579306 -340 579374 -284
rect 579430 -340 579498 -284
rect 579554 -340 579622 -284
rect 579678 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect -956 -408 597020 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 3250 -408
rect 3306 -464 3374 -408
rect 3430 -464 3498 -408
rect 3554 -464 3622 -408
rect 3678 -464 21250 -408
rect 21306 -464 21374 -408
rect 21430 -464 21498 -408
rect 21554 -464 21622 -408
rect 21678 -464 39250 -408
rect 39306 -464 39374 -408
rect 39430 -464 39498 -408
rect 39554 -464 39622 -408
rect 39678 -464 57250 -408
rect 57306 -464 57374 -408
rect 57430 -464 57498 -408
rect 57554 -464 57622 -408
rect 57678 -464 75250 -408
rect 75306 -464 75374 -408
rect 75430 -464 75498 -408
rect 75554 -464 75622 -408
rect 75678 -464 93250 -408
rect 93306 -464 93374 -408
rect 93430 -464 93498 -408
rect 93554 -464 93622 -408
rect 93678 -464 111250 -408
rect 111306 -464 111374 -408
rect 111430 -464 111498 -408
rect 111554 -464 111622 -408
rect 111678 -464 129250 -408
rect 129306 -464 129374 -408
rect 129430 -464 129498 -408
rect 129554 -464 129622 -408
rect 129678 -464 147250 -408
rect 147306 -464 147374 -408
rect 147430 -464 147498 -408
rect 147554 -464 147622 -408
rect 147678 -464 165250 -408
rect 165306 -464 165374 -408
rect 165430 -464 165498 -408
rect 165554 -464 165622 -408
rect 165678 -464 183250 -408
rect 183306 -464 183374 -408
rect 183430 -464 183498 -408
rect 183554 -464 183622 -408
rect 183678 -464 201250 -408
rect 201306 -464 201374 -408
rect 201430 -464 201498 -408
rect 201554 -464 201622 -408
rect 201678 -464 219250 -408
rect 219306 -464 219374 -408
rect 219430 -464 219498 -408
rect 219554 -464 219622 -408
rect 219678 -464 237250 -408
rect 237306 -464 237374 -408
rect 237430 -464 237498 -408
rect 237554 -464 237622 -408
rect 237678 -464 255250 -408
rect 255306 -464 255374 -408
rect 255430 -464 255498 -408
rect 255554 -464 255622 -408
rect 255678 -464 273250 -408
rect 273306 -464 273374 -408
rect 273430 -464 273498 -408
rect 273554 -464 273622 -408
rect 273678 -464 291250 -408
rect 291306 -464 291374 -408
rect 291430 -464 291498 -408
rect 291554 -464 291622 -408
rect 291678 -464 309250 -408
rect 309306 -464 309374 -408
rect 309430 -464 309498 -408
rect 309554 -464 309622 -408
rect 309678 -464 327250 -408
rect 327306 -464 327374 -408
rect 327430 -464 327498 -408
rect 327554 -464 327622 -408
rect 327678 -464 345250 -408
rect 345306 -464 345374 -408
rect 345430 -464 345498 -408
rect 345554 -464 345622 -408
rect 345678 -464 363250 -408
rect 363306 -464 363374 -408
rect 363430 -464 363498 -408
rect 363554 -464 363622 -408
rect 363678 -464 381250 -408
rect 381306 -464 381374 -408
rect 381430 -464 381498 -408
rect 381554 -464 381622 -408
rect 381678 -464 399250 -408
rect 399306 -464 399374 -408
rect 399430 -464 399498 -408
rect 399554 -464 399622 -408
rect 399678 -464 417250 -408
rect 417306 -464 417374 -408
rect 417430 -464 417498 -408
rect 417554 -464 417622 -408
rect 417678 -464 435250 -408
rect 435306 -464 435374 -408
rect 435430 -464 435498 -408
rect 435554 -464 435622 -408
rect 435678 -464 453250 -408
rect 453306 -464 453374 -408
rect 453430 -464 453498 -408
rect 453554 -464 453622 -408
rect 453678 -464 471250 -408
rect 471306 -464 471374 -408
rect 471430 -464 471498 -408
rect 471554 -464 471622 -408
rect 471678 -464 489250 -408
rect 489306 -464 489374 -408
rect 489430 -464 489498 -408
rect 489554 -464 489622 -408
rect 489678 -464 507250 -408
rect 507306 -464 507374 -408
rect 507430 -464 507498 -408
rect 507554 -464 507622 -408
rect 507678 -464 525250 -408
rect 525306 -464 525374 -408
rect 525430 -464 525498 -408
rect 525554 -464 525622 -408
rect 525678 -464 543250 -408
rect 543306 -464 543374 -408
rect 543430 -464 543498 -408
rect 543554 -464 543622 -408
rect 543678 -464 561250 -408
rect 561306 -464 561374 -408
rect 561430 -464 561498 -408
rect 561554 -464 561622 -408
rect 561678 -464 579250 -408
rect 579306 -464 579374 -408
rect 579430 -464 579498 -408
rect 579554 -464 579622 -408
rect 579678 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect -956 -532 597020 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 3250 -532
rect 3306 -588 3374 -532
rect 3430 -588 3498 -532
rect 3554 -588 3622 -532
rect 3678 -588 21250 -532
rect 21306 -588 21374 -532
rect 21430 -588 21498 -532
rect 21554 -588 21622 -532
rect 21678 -588 39250 -532
rect 39306 -588 39374 -532
rect 39430 -588 39498 -532
rect 39554 -588 39622 -532
rect 39678 -588 57250 -532
rect 57306 -588 57374 -532
rect 57430 -588 57498 -532
rect 57554 -588 57622 -532
rect 57678 -588 75250 -532
rect 75306 -588 75374 -532
rect 75430 -588 75498 -532
rect 75554 -588 75622 -532
rect 75678 -588 93250 -532
rect 93306 -588 93374 -532
rect 93430 -588 93498 -532
rect 93554 -588 93622 -532
rect 93678 -588 111250 -532
rect 111306 -588 111374 -532
rect 111430 -588 111498 -532
rect 111554 -588 111622 -532
rect 111678 -588 129250 -532
rect 129306 -588 129374 -532
rect 129430 -588 129498 -532
rect 129554 -588 129622 -532
rect 129678 -588 147250 -532
rect 147306 -588 147374 -532
rect 147430 -588 147498 -532
rect 147554 -588 147622 -532
rect 147678 -588 165250 -532
rect 165306 -588 165374 -532
rect 165430 -588 165498 -532
rect 165554 -588 165622 -532
rect 165678 -588 183250 -532
rect 183306 -588 183374 -532
rect 183430 -588 183498 -532
rect 183554 -588 183622 -532
rect 183678 -588 201250 -532
rect 201306 -588 201374 -532
rect 201430 -588 201498 -532
rect 201554 -588 201622 -532
rect 201678 -588 219250 -532
rect 219306 -588 219374 -532
rect 219430 -588 219498 -532
rect 219554 -588 219622 -532
rect 219678 -588 237250 -532
rect 237306 -588 237374 -532
rect 237430 -588 237498 -532
rect 237554 -588 237622 -532
rect 237678 -588 255250 -532
rect 255306 -588 255374 -532
rect 255430 -588 255498 -532
rect 255554 -588 255622 -532
rect 255678 -588 273250 -532
rect 273306 -588 273374 -532
rect 273430 -588 273498 -532
rect 273554 -588 273622 -532
rect 273678 -588 291250 -532
rect 291306 -588 291374 -532
rect 291430 -588 291498 -532
rect 291554 -588 291622 -532
rect 291678 -588 309250 -532
rect 309306 -588 309374 -532
rect 309430 -588 309498 -532
rect 309554 -588 309622 -532
rect 309678 -588 327250 -532
rect 327306 -588 327374 -532
rect 327430 -588 327498 -532
rect 327554 -588 327622 -532
rect 327678 -588 345250 -532
rect 345306 -588 345374 -532
rect 345430 -588 345498 -532
rect 345554 -588 345622 -532
rect 345678 -588 363250 -532
rect 363306 -588 363374 -532
rect 363430 -588 363498 -532
rect 363554 -588 363622 -532
rect 363678 -588 381250 -532
rect 381306 -588 381374 -532
rect 381430 -588 381498 -532
rect 381554 -588 381622 -532
rect 381678 -588 399250 -532
rect 399306 -588 399374 -532
rect 399430 -588 399498 -532
rect 399554 -588 399622 -532
rect 399678 -588 417250 -532
rect 417306 -588 417374 -532
rect 417430 -588 417498 -532
rect 417554 -588 417622 -532
rect 417678 -588 435250 -532
rect 435306 -588 435374 -532
rect 435430 -588 435498 -532
rect 435554 -588 435622 -532
rect 435678 -588 453250 -532
rect 453306 -588 453374 -532
rect 453430 -588 453498 -532
rect 453554 -588 453622 -532
rect 453678 -588 471250 -532
rect 471306 -588 471374 -532
rect 471430 -588 471498 -532
rect 471554 -588 471622 -532
rect 471678 -588 489250 -532
rect 489306 -588 489374 -532
rect 489430 -588 489498 -532
rect 489554 -588 489622 -532
rect 489678 -588 507250 -532
rect 507306 -588 507374 -532
rect 507430 -588 507498 -532
rect 507554 -588 507622 -532
rect 507678 -588 525250 -532
rect 525306 -588 525374 -532
rect 525430 -588 525498 -532
rect 525554 -588 525622 -532
rect 525678 -588 543250 -532
rect 543306 -588 543374 -532
rect 543430 -588 543498 -532
rect 543554 -588 543622 -532
rect 543678 -588 561250 -532
rect 561306 -588 561374 -532
rect 561430 -588 561498 -532
rect 561554 -588 561622 -532
rect 561678 -588 579250 -532
rect 579306 -588 579374 -532
rect 579430 -588 579498 -532
rect 579554 -588 579622 -532
rect 579678 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect -956 -684 597020 -588
rect -1916 -1120 597980 -1024
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 6970 -1120
rect 7026 -1176 7094 -1120
rect 7150 -1176 7218 -1120
rect 7274 -1176 7342 -1120
rect 7398 -1176 24970 -1120
rect 25026 -1176 25094 -1120
rect 25150 -1176 25218 -1120
rect 25274 -1176 25342 -1120
rect 25398 -1176 42970 -1120
rect 43026 -1176 43094 -1120
rect 43150 -1176 43218 -1120
rect 43274 -1176 43342 -1120
rect 43398 -1176 60970 -1120
rect 61026 -1176 61094 -1120
rect 61150 -1176 61218 -1120
rect 61274 -1176 61342 -1120
rect 61398 -1176 78970 -1120
rect 79026 -1176 79094 -1120
rect 79150 -1176 79218 -1120
rect 79274 -1176 79342 -1120
rect 79398 -1176 96970 -1120
rect 97026 -1176 97094 -1120
rect 97150 -1176 97218 -1120
rect 97274 -1176 97342 -1120
rect 97398 -1176 114970 -1120
rect 115026 -1176 115094 -1120
rect 115150 -1176 115218 -1120
rect 115274 -1176 115342 -1120
rect 115398 -1176 132970 -1120
rect 133026 -1176 133094 -1120
rect 133150 -1176 133218 -1120
rect 133274 -1176 133342 -1120
rect 133398 -1176 150970 -1120
rect 151026 -1176 151094 -1120
rect 151150 -1176 151218 -1120
rect 151274 -1176 151342 -1120
rect 151398 -1176 168970 -1120
rect 169026 -1176 169094 -1120
rect 169150 -1176 169218 -1120
rect 169274 -1176 169342 -1120
rect 169398 -1176 186970 -1120
rect 187026 -1176 187094 -1120
rect 187150 -1176 187218 -1120
rect 187274 -1176 187342 -1120
rect 187398 -1176 204970 -1120
rect 205026 -1176 205094 -1120
rect 205150 -1176 205218 -1120
rect 205274 -1176 205342 -1120
rect 205398 -1176 222970 -1120
rect 223026 -1176 223094 -1120
rect 223150 -1176 223218 -1120
rect 223274 -1176 223342 -1120
rect 223398 -1176 240970 -1120
rect 241026 -1176 241094 -1120
rect 241150 -1176 241218 -1120
rect 241274 -1176 241342 -1120
rect 241398 -1176 258970 -1120
rect 259026 -1176 259094 -1120
rect 259150 -1176 259218 -1120
rect 259274 -1176 259342 -1120
rect 259398 -1176 276970 -1120
rect 277026 -1176 277094 -1120
rect 277150 -1176 277218 -1120
rect 277274 -1176 277342 -1120
rect 277398 -1176 294970 -1120
rect 295026 -1176 295094 -1120
rect 295150 -1176 295218 -1120
rect 295274 -1176 295342 -1120
rect 295398 -1176 312970 -1120
rect 313026 -1176 313094 -1120
rect 313150 -1176 313218 -1120
rect 313274 -1176 313342 -1120
rect 313398 -1176 330970 -1120
rect 331026 -1176 331094 -1120
rect 331150 -1176 331218 -1120
rect 331274 -1176 331342 -1120
rect 331398 -1176 348970 -1120
rect 349026 -1176 349094 -1120
rect 349150 -1176 349218 -1120
rect 349274 -1176 349342 -1120
rect 349398 -1176 366970 -1120
rect 367026 -1176 367094 -1120
rect 367150 -1176 367218 -1120
rect 367274 -1176 367342 -1120
rect 367398 -1176 384970 -1120
rect 385026 -1176 385094 -1120
rect 385150 -1176 385218 -1120
rect 385274 -1176 385342 -1120
rect 385398 -1176 402970 -1120
rect 403026 -1176 403094 -1120
rect 403150 -1176 403218 -1120
rect 403274 -1176 403342 -1120
rect 403398 -1176 420970 -1120
rect 421026 -1176 421094 -1120
rect 421150 -1176 421218 -1120
rect 421274 -1176 421342 -1120
rect 421398 -1176 438970 -1120
rect 439026 -1176 439094 -1120
rect 439150 -1176 439218 -1120
rect 439274 -1176 439342 -1120
rect 439398 -1176 456970 -1120
rect 457026 -1176 457094 -1120
rect 457150 -1176 457218 -1120
rect 457274 -1176 457342 -1120
rect 457398 -1176 474970 -1120
rect 475026 -1176 475094 -1120
rect 475150 -1176 475218 -1120
rect 475274 -1176 475342 -1120
rect 475398 -1176 492970 -1120
rect 493026 -1176 493094 -1120
rect 493150 -1176 493218 -1120
rect 493274 -1176 493342 -1120
rect 493398 -1176 510970 -1120
rect 511026 -1176 511094 -1120
rect 511150 -1176 511218 -1120
rect 511274 -1176 511342 -1120
rect 511398 -1176 528970 -1120
rect 529026 -1176 529094 -1120
rect 529150 -1176 529218 -1120
rect 529274 -1176 529342 -1120
rect 529398 -1176 546970 -1120
rect 547026 -1176 547094 -1120
rect 547150 -1176 547218 -1120
rect 547274 -1176 547342 -1120
rect 547398 -1176 564970 -1120
rect 565026 -1176 565094 -1120
rect 565150 -1176 565218 -1120
rect 565274 -1176 565342 -1120
rect 565398 -1176 582970 -1120
rect 583026 -1176 583094 -1120
rect 583150 -1176 583218 -1120
rect 583274 -1176 583342 -1120
rect 583398 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect -1916 -1244 597980 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 6970 -1244
rect 7026 -1300 7094 -1244
rect 7150 -1300 7218 -1244
rect 7274 -1300 7342 -1244
rect 7398 -1300 24970 -1244
rect 25026 -1300 25094 -1244
rect 25150 -1300 25218 -1244
rect 25274 -1300 25342 -1244
rect 25398 -1300 42970 -1244
rect 43026 -1300 43094 -1244
rect 43150 -1300 43218 -1244
rect 43274 -1300 43342 -1244
rect 43398 -1300 60970 -1244
rect 61026 -1300 61094 -1244
rect 61150 -1300 61218 -1244
rect 61274 -1300 61342 -1244
rect 61398 -1300 78970 -1244
rect 79026 -1300 79094 -1244
rect 79150 -1300 79218 -1244
rect 79274 -1300 79342 -1244
rect 79398 -1300 96970 -1244
rect 97026 -1300 97094 -1244
rect 97150 -1300 97218 -1244
rect 97274 -1300 97342 -1244
rect 97398 -1300 114970 -1244
rect 115026 -1300 115094 -1244
rect 115150 -1300 115218 -1244
rect 115274 -1300 115342 -1244
rect 115398 -1300 132970 -1244
rect 133026 -1300 133094 -1244
rect 133150 -1300 133218 -1244
rect 133274 -1300 133342 -1244
rect 133398 -1300 150970 -1244
rect 151026 -1300 151094 -1244
rect 151150 -1300 151218 -1244
rect 151274 -1300 151342 -1244
rect 151398 -1300 168970 -1244
rect 169026 -1300 169094 -1244
rect 169150 -1300 169218 -1244
rect 169274 -1300 169342 -1244
rect 169398 -1300 186970 -1244
rect 187026 -1300 187094 -1244
rect 187150 -1300 187218 -1244
rect 187274 -1300 187342 -1244
rect 187398 -1300 204970 -1244
rect 205026 -1300 205094 -1244
rect 205150 -1300 205218 -1244
rect 205274 -1300 205342 -1244
rect 205398 -1300 222970 -1244
rect 223026 -1300 223094 -1244
rect 223150 -1300 223218 -1244
rect 223274 -1300 223342 -1244
rect 223398 -1300 240970 -1244
rect 241026 -1300 241094 -1244
rect 241150 -1300 241218 -1244
rect 241274 -1300 241342 -1244
rect 241398 -1300 258970 -1244
rect 259026 -1300 259094 -1244
rect 259150 -1300 259218 -1244
rect 259274 -1300 259342 -1244
rect 259398 -1300 276970 -1244
rect 277026 -1300 277094 -1244
rect 277150 -1300 277218 -1244
rect 277274 -1300 277342 -1244
rect 277398 -1300 294970 -1244
rect 295026 -1300 295094 -1244
rect 295150 -1300 295218 -1244
rect 295274 -1300 295342 -1244
rect 295398 -1300 312970 -1244
rect 313026 -1300 313094 -1244
rect 313150 -1300 313218 -1244
rect 313274 -1300 313342 -1244
rect 313398 -1300 330970 -1244
rect 331026 -1300 331094 -1244
rect 331150 -1300 331218 -1244
rect 331274 -1300 331342 -1244
rect 331398 -1300 348970 -1244
rect 349026 -1300 349094 -1244
rect 349150 -1300 349218 -1244
rect 349274 -1300 349342 -1244
rect 349398 -1300 366970 -1244
rect 367026 -1300 367094 -1244
rect 367150 -1300 367218 -1244
rect 367274 -1300 367342 -1244
rect 367398 -1300 384970 -1244
rect 385026 -1300 385094 -1244
rect 385150 -1300 385218 -1244
rect 385274 -1300 385342 -1244
rect 385398 -1300 402970 -1244
rect 403026 -1300 403094 -1244
rect 403150 -1300 403218 -1244
rect 403274 -1300 403342 -1244
rect 403398 -1300 420970 -1244
rect 421026 -1300 421094 -1244
rect 421150 -1300 421218 -1244
rect 421274 -1300 421342 -1244
rect 421398 -1300 438970 -1244
rect 439026 -1300 439094 -1244
rect 439150 -1300 439218 -1244
rect 439274 -1300 439342 -1244
rect 439398 -1300 456970 -1244
rect 457026 -1300 457094 -1244
rect 457150 -1300 457218 -1244
rect 457274 -1300 457342 -1244
rect 457398 -1300 474970 -1244
rect 475026 -1300 475094 -1244
rect 475150 -1300 475218 -1244
rect 475274 -1300 475342 -1244
rect 475398 -1300 492970 -1244
rect 493026 -1300 493094 -1244
rect 493150 -1300 493218 -1244
rect 493274 -1300 493342 -1244
rect 493398 -1300 510970 -1244
rect 511026 -1300 511094 -1244
rect 511150 -1300 511218 -1244
rect 511274 -1300 511342 -1244
rect 511398 -1300 528970 -1244
rect 529026 -1300 529094 -1244
rect 529150 -1300 529218 -1244
rect 529274 -1300 529342 -1244
rect 529398 -1300 546970 -1244
rect 547026 -1300 547094 -1244
rect 547150 -1300 547218 -1244
rect 547274 -1300 547342 -1244
rect 547398 -1300 564970 -1244
rect 565026 -1300 565094 -1244
rect 565150 -1300 565218 -1244
rect 565274 -1300 565342 -1244
rect 565398 -1300 582970 -1244
rect 583026 -1300 583094 -1244
rect 583150 -1300 583218 -1244
rect 583274 -1300 583342 -1244
rect 583398 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect -1916 -1368 597980 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 6970 -1368
rect 7026 -1424 7094 -1368
rect 7150 -1424 7218 -1368
rect 7274 -1424 7342 -1368
rect 7398 -1424 24970 -1368
rect 25026 -1424 25094 -1368
rect 25150 -1424 25218 -1368
rect 25274 -1424 25342 -1368
rect 25398 -1424 42970 -1368
rect 43026 -1424 43094 -1368
rect 43150 -1424 43218 -1368
rect 43274 -1424 43342 -1368
rect 43398 -1424 60970 -1368
rect 61026 -1424 61094 -1368
rect 61150 -1424 61218 -1368
rect 61274 -1424 61342 -1368
rect 61398 -1424 78970 -1368
rect 79026 -1424 79094 -1368
rect 79150 -1424 79218 -1368
rect 79274 -1424 79342 -1368
rect 79398 -1424 96970 -1368
rect 97026 -1424 97094 -1368
rect 97150 -1424 97218 -1368
rect 97274 -1424 97342 -1368
rect 97398 -1424 114970 -1368
rect 115026 -1424 115094 -1368
rect 115150 -1424 115218 -1368
rect 115274 -1424 115342 -1368
rect 115398 -1424 132970 -1368
rect 133026 -1424 133094 -1368
rect 133150 -1424 133218 -1368
rect 133274 -1424 133342 -1368
rect 133398 -1424 150970 -1368
rect 151026 -1424 151094 -1368
rect 151150 -1424 151218 -1368
rect 151274 -1424 151342 -1368
rect 151398 -1424 168970 -1368
rect 169026 -1424 169094 -1368
rect 169150 -1424 169218 -1368
rect 169274 -1424 169342 -1368
rect 169398 -1424 186970 -1368
rect 187026 -1424 187094 -1368
rect 187150 -1424 187218 -1368
rect 187274 -1424 187342 -1368
rect 187398 -1424 204970 -1368
rect 205026 -1424 205094 -1368
rect 205150 -1424 205218 -1368
rect 205274 -1424 205342 -1368
rect 205398 -1424 222970 -1368
rect 223026 -1424 223094 -1368
rect 223150 -1424 223218 -1368
rect 223274 -1424 223342 -1368
rect 223398 -1424 240970 -1368
rect 241026 -1424 241094 -1368
rect 241150 -1424 241218 -1368
rect 241274 -1424 241342 -1368
rect 241398 -1424 258970 -1368
rect 259026 -1424 259094 -1368
rect 259150 -1424 259218 -1368
rect 259274 -1424 259342 -1368
rect 259398 -1424 276970 -1368
rect 277026 -1424 277094 -1368
rect 277150 -1424 277218 -1368
rect 277274 -1424 277342 -1368
rect 277398 -1424 294970 -1368
rect 295026 -1424 295094 -1368
rect 295150 -1424 295218 -1368
rect 295274 -1424 295342 -1368
rect 295398 -1424 312970 -1368
rect 313026 -1424 313094 -1368
rect 313150 -1424 313218 -1368
rect 313274 -1424 313342 -1368
rect 313398 -1424 330970 -1368
rect 331026 -1424 331094 -1368
rect 331150 -1424 331218 -1368
rect 331274 -1424 331342 -1368
rect 331398 -1424 348970 -1368
rect 349026 -1424 349094 -1368
rect 349150 -1424 349218 -1368
rect 349274 -1424 349342 -1368
rect 349398 -1424 366970 -1368
rect 367026 -1424 367094 -1368
rect 367150 -1424 367218 -1368
rect 367274 -1424 367342 -1368
rect 367398 -1424 384970 -1368
rect 385026 -1424 385094 -1368
rect 385150 -1424 385218 -1368
rect 385274 -1424 385342 -1368
rect 385398 -1424 402970 -1368
rect 403026 -1424 403094 -1368
rect 403150 -1424 403218 -1368
rect 403274 -1424 403342 -1368
rect 403398 -1424 420970 -1368
rect 421026 -1424 421094 -1368
rect 421150 -1424 421218 -1368
rect 421274 -1424 421342 -1368
rect 421398 -1424 438970 -1368
rect 439026 -1424 439094 -1368
rect 439150 -1424 439218 -1368
rect 439274 -1424 439342 -1368
rect 439398 -1424 456970 -1368
rect 457026 -1424 457094 -1368
rect 457150 -1424 457218 -1368
rect 457274 -1424 457342 -1368
rect 457398 -1424 474970 -1368
rect 475026 -1424 475094 -1368
rect 475150 -1424 475218 -1368
rect 475274 -1424 475342 -1368
rect 475398 -1424 492970 -1368
rect 493026 -1424 493094 -1368
rect 493150 -1424 493218 -1368
rect 493274 -1424 493342 -1368
rect 493398 -1424 510970 -1368
rect 511026 -1424 511094 -1368
rect 511150 -1424 511218 -1368
rect 511274 -1424 511342 -1368
rect 511398 -1424 528970 -1368
rect 529026 -1424 529094 -1368
rect 529150 -1424 529218 -1368
rect 529274 -1424 529342 -1368
rect 529398 -1424 546970 -1368
rect 547026 -1424 547094 -1368
rect 547150 -1424 547218 -1368
rect 547274 -1424 547342 -1368
rect 547398 -1424 564970 -1368
rect 565026 -1424 565094 -1368
rect 565150 -1424 565218 -1368
rect 565274 -1424 565342 -1368
rect 565398 -1424 582970 -1368
rect 583026 -1424 583094 -1368
rect 583150 -1424 583218 -1368
rect 583274 -1424 583342 -1368
rect 583398 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect -1916 -1492 597980 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 6970 -1492
rect 7026 -1548 7094 -1492
rect 7150 -1548 7218 -1492
rect 7274 -1548 7342 -1492
rect 7398 -1548 24970 -1492
rect 25026 -1548 25094 -1492
rect 25150 -1548 25218 -1492
rect 25274 -1548 25342 -1492
rect 25398 -1548 42970 -1492
rect 43026 -1548 43094 -1492
rect 43150 -1548 43218 -1492
rect 43274 -1548 43342 -1492
rect 43398 -1548 60970 -1492
rect 61026 -1548 61094 -1492
rect 61150 -1548 61218 -1492
rect 61274 -1548 61342 -1492
rect 61398 -1548 78970 -1492
rect 79026 -1548 79094 -1492
rect 79150 -1548 79218 -1492
rect 79274 -1548 79342 -1492
rect 79398 -1548 96970 -1492
rect 97026 -1548 97094 -1492
rect 97150 -1548 97218 -1492
rect 97274 -1548 97342 -1492
rect 97398 -1548 114970 -1492
rect 115026 -1548 115094 -1492
rect 115150 -1548 115218 -1492
rect 115274 -1548 115342 -1492
rect 115398 -1548 132970 -1492
rect 133026 -1548 133094 -1492
rect 133150 -1548 133218 -1492
rect 133274 -1548 133342 -1492
rect 133398 -1548 150970 -1492
rect 151026 -1548 151094 -1492
rect 151150 -1548 151218 -1492
rect 151274 -1548 151342 -1492
rect 151398 -1548 168970 -1492
rect 169026 -1548 169094 -1492
rect 169150 -1548 169218 -1492
rect 169274 -1548 169342 -1492
rect 169398 -1548 186970 -1492
rect 187026 -1548 187094 -1492
rect 187150 -1548 187218 -1492
rect 187274 -1548 187342 -1492
rect 187398 -1548 204970 -1492
rect 205026 -1548 205094 -1492
rect 205150 -1548 205218 -1492
rect 205274 -1548 205342 -1492
rect 205398 -1548 222970 -1492
rect 223026 -1548 223094 -1492
rect 223150 -1548 223218 -1492
rect 223274 -1548 223342 -1492
rect 223398 -1548 240970 -1492
rect 241026 -1548 241094 -1492
rect 241150 -1548 241218 -1492
rect 241274 -1548 241342 -1492
rect 241398 -1548 258970 -1492
rect 259026 -1548 259094 -1492
rect 259150 -1548 259218 -1492
rect 259274 -1548 259342 -1492
rect 259398 -1548 276970 -1492
rect 277026 -1548 277094 -1492
rect 277150 -1548 277218 -1492
rect 277274 -1548 277342 -1492
rect 277398 -1548 294970 -1492
rect 295026 -1548 295094 -1492
rect 295150 -1548 295218 -1492
rect 295274 -1548 295342 -1492
rect 295398 -1548 312970 -1492
rect 313026 -1548 313094 -1492
rect 313150 -1548 313218 -1492
rect 313274 -1548 313342 -1492
rect 313398 -1548 330970 -1492
rect 331026 -1548 331094 -1492
rect 331150 -1548 331218 -1492
rect 331274 -1548 331342 -1492
rect 331398 -1548 348970 -1492
rect 349026 -1548 349094 -1492
rect 349150 -1548 349218 -1492
rect 349274 -1548 349342 -1492
rect 349398 -1548 366970 -1492
rect 367026 -1548 367094 -1492
rect 367150 -1548 367218 -1492
rect 367274 -1548 367342 -1492
rect 367398 -1548 384970 -1492
rect 385026 -1548 385094 -1492
rect 385150 -1548 385218 -1492
rect 385274 -1548 385342 -1492
rect 385398 -1548 402970 -1492
rect 403026 -1548 403094 -1492
rect 403150 -1548 403218 -1492
rect 403274 -1548 403342 -1492
rect 403398 -1548 420970 -1492
rect 421026 -1548 421094 -1492
rect 421150 -1548 421218 -1492
rect 421274 -1548 421342 -1492
rect 421398 -1548 438970 -1492
rect 439026 -1548 439094 -1492
rect 439150 -1548 439218 -1492
rect 439274 -1548 439342 -1492
rect 439398 -1548 456970 -1492
rect 457026 -1548 457094 -1492
rect 457150 -1548 457218 -1492
rect 457274 -1548 457342 -1492
rect 457398 -1548 474970 -1492
rect 475026 -1548 475094 -1492
rect 475150 -1548 475218 -1492
rect 475274 -1548 475342 -1492
rect 475398 -1548 492970 -1492
rect 493026 -1548 493094 -1492
rect 493150 -1548 493218 -1492
rect 493274 -1548 493342 -1492
rect 493398 -1548 510970 -1492
rect 511026 -1548 511094 -1492
rect 511150 -1548 511218 -1492
rect 511274 -1548 511342 -1492
rect 511398 -1548 528970 -1492
rect 529026 -1548 529094 -1492
rect 529150 -1548 529218 -1492
rect 529274 -1548 529342 -1492
rect 529398 -1548 546970 -1492
rect 547026 -1548 547094 -1492
rect 547150 -1548 547218 -1492
rect 547274 -1548 547342 -1492
rect 547398 -1548 564970 -1492
rect 565026 -1548 565094 -1492
rect 565150 -1548 565218 -1492
rect 565274 -1548 565342 -1492
rect 565398 -1548 582970 -1492
rect 583026 -1548 583094 -1492
rect 583150 -1548 583218 -1492
rect 583274 -1548 583342 -1492
rect 583398 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect -1916 -1644 597980 -1548
use aes128  aes128
timestamp 0
transform 1 0 50000 0 1 30000
box 0 200 499940 499940
<< labels >>
flabel metal3 s 595560 7112 597000 7336 0 FreeSans 896 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 595560 403592 597000 403816 0 FreeSans 896 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 595560 443240 597000 443464 0 FreeSans 896 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 595560 482888 597000 483112 0 FreeSans 896 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 595560 522536 597000 522760 0 FreeSans 896 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 595560 562184 597000 562408 0 FreeSans 896 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 584696 595560 584920 597000 0 FreeSans 896 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 518504 595560 518728 597000 0 FreeSans 896 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 452312 595560 452536 597000 0 FreeSans 896 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 386120 595560 386344 597000 0 FreeSans 896 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 319928 595560 320152 597000 0 FreeSans 896 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 595560 46760 597000 46984 0 FreeSans 896 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 253736 595560 253960 597000 0 FreeSans 896 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 187544 595560 187768 597000 0 FreeSans 896 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 121352 595560 121576 597000 0 FreeSans 896 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 55160 595560 55384 597000 0 FreeSans 896 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s -960 587160 480 587384 0 FreeSans 896 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s -960 544824 480 545048 0 FreeSans 896 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s -960 502488 480 502712 0 FreeSans 896 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s -960 460152 480 460376 0 FreeSans 896 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s -960 417816 480 418040 0 FreeSans 896 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s -960 375480 480 375704 0 FreeSans 896 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 595560 86408 597000 86632 0 FreeSans 896 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s -960 333144 480 333368 0 FreeSans 896 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s -960 290808 480 291032 0 FreeSans 896 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s -960 248472 480 248696 0 FreeSans 896 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s -960 206136 480 206360 0 FreeSans 896 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s -960 163800 480 164024 0 FreeSans 896 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s -960 121464 480 121688 0 FreeSans 896 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s -960 79128 480 79352 0 FreeSans 896 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s -960 36792 480 37016 0 FreeSans 896 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 595560 126056 597000 126280 0 FreeSans 896 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 595560 165704 597000 165928 0 FreeSans 896 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 595560 205352 597000 205576 0 FreeSans 896 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 595560 245000 597000 245224 0 FreeSans 896 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 595560 284648 597000 284872 0 FreeSans 896 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 595560 324296 597000 324520 0 FreeSans 896 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 595560 363944 597000 364168 0 FreeSans 896 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal3 s 595560 33544 597000 33768 0 FreeSans 896 0 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 595560 430024 597000 430248 0 FreeSans 896 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 595560 469672 597000 469896 0 FreeSans 896 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 595560 509320 597000 509544 0 FreeSans 896 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 595560 548968 597000 549192 0 FreeSans 896 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 595560 588616 597000 588840 0 FreeSans 896 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 540568 595560 540792 597000 0 FreeSans 896 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 474376 595560 474600 597000 0 FreeSans 896 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 408184 595560 408408 597000 0 FreeSans 896 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 341992 595560 342216 597000 0 FreeSans 896 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 275800 595560 276024 597000 0 FreeSans 896 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal3 s 595560 73192 597000 73416 0 FreeSans 896 0 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 209608 595560 209832 597000 0 FreeSans 896 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 143416 595560 143640 597000 0 FreeSans 896 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 77224 595560 77448 597000 0 FreeSans 896 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 11032 595560 11256 597000 0 FreeSans 896 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s -960 558936 480 559160 0 FreeSans 896 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal3 s -960 516600 480 516824 0 FreeSans 896 0 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal3 s -960 474264 480 474488 0 FreeSans 896 0 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s -960 431928 480 432152 0 FreeSans 896 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s -960 389592 480 389816 0 FreeSans 896 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s -960 347256 480 347480 0 FreeSans 896 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal3 s 595560 112840 597000 113064 0 FreeSans 896 0 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal3 s -960 304920 480 305144 0 FreeSans 896 0 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s -960 262584 480 262808 0 FreeSans 896 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s -960 220248 480 220472 0 FreeSans 896 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s -960 177912 480 178136 0 FreeSans 896 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s -960 135576 480 135800 0 FreeSans 896 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s -960 93240 480 93464 0 FreeSans 896 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal3 s -960 50904 480 51128 0 FreeSans 896 0 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s -960 8568 480 8792 0 FreeSans 896 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 595560 152488 597000 152712 0 FreeSans 896 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal3 s 595560 192136 597000 192360 0 FreeSans 896 0 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 595560 231784 597000 232008 0 FreeSans 896 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 595560 271432 597000 271656 0 FreeSans 896 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 595560 311080 597000 311304 0 FreeSans 896 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 595560 350728 597000 350952 0 FreeSans 896 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal3 s 595560 390376 597000 390600 0 FreeSans 896 0 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 595560 20328 597000 20552 0 FreeSans 896 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 595560 416808 597000 417032 0 FreeSans 896 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 595560 456456 597000 456680 0 FreeSans 896 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 595560 496104 597000 496328 0 FreeSans 896 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 595560 535752 597000 535976 0 FreeSans 896 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal3 s 595560 575400 597000 575624 0 FreeSans 896 0 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 562632 595560 562856 597000 0 FreeSans 896 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 496440 595560 496664 597000 0 FreeSans 896 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 430248 595560 430472 597000 0 FreeSans 896 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 364056 595560 364280 597000 0 FreeSans 896 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 297864 595560 298088 597000 0 FreeSans 896 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal3 s 595560 59976 597000 60200 0 FreeSans 896 0 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 231672 595560 231896 597000 0 FreeSans 896 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 165480 595560 165704 597000 0 FreeSans 896 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 99288 595560 99512 597000 0 FreeSans 896 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 33096 595560 33320 597000 0 FreeSans 896 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s -960 573048 480 573272 0 FreeSans 896 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal3 s -960 530712 480 530936 0 FreeSans 896 0 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal3 s -960 488376 480 488600 0 FreeSans 896 0 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal3 s -960 446040 480 446264 0 FreeSans 896 0 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal3 s -960 403704 480 403928 0 FreeSans 896 0 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal3 s -960 361368 480 361592 0 FreeSans 896 0 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 595560 99624 597000 99848 0 FreeSans 896 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s -960 319032 480 319256 0 FreeSans 896 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s -960 276696 480 276920 0 FreeSans 896 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal3 s -960 234360 480 234584 0 FreeSans 896 0 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal3 s -960 192024 480 192248 0 FreeSans 896 0 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s -960 149688 480 149912 0 FreeSans 896 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s -960 107352 480 107576 0 FreeSans 896 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal3 s -960 65016 480 65240 0 FreeSans 896 0 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s -960 22680 480 22904 0 FreeSans 896 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal3 s 595560 139272 597000 139496 0 FreeSans 896 0 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal3 s 595560 178920 597000 179144 0 FreeSans 896 0 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal3 s 595560 218568 597000 218792 0 FreeSans 896 0 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 595560 258216 597000 258440 0 FreeSans 896 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 595560 297864 597000 298088 0 FreeSans 896 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 595560 337512 597000 337736 0 FreeSans 896 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 595560 377160 597000 377384 0 FreeSans 896 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal2 s 213192 -960 213416 480 0 FreeSans 896 90 0 0 la_data_in[0]
port 114 nsew signal input
flabel metal2 s 270312 -960 270536 480 0 FreeSans 896 90 0 0 la_data_in[10]
port 115 nsew signal input
flabel metal2 s 276024 -960 276248 480 0 FreeSans 896 90 0 0 la_data_in[11]
port 116 nsew signal input
flabel metal2 s 281736 -960 281960 480 0 FreeSans 896 90 0 0 la_data_in[12]
port 117 nsew signal input
flabel metal2 s 287448 -960 287672 480 0 FreeSans 896 90 0 0 la_data_in[13]
port 118 nsew signal input
flabel metal2 s 293160 -960 293384 480 0 FreeSans 896 90 0 0 la_data_in[14]
port 119 nsew signal input
flabel metal2 s 298872 -960 299096 480 0 FreeSans 896 90 0 0 la_data_in[15]
port 120 nsew signal input
flabel metal2 s 304584 -960 304808 480 0 FreeSans 896 90 0 0 la_data_in[16]
port 121 nsew signal input
flabel metal2 s 310296 -960 310520 480 0 FreeSans 896 90 0 0 la_data_in[17]
port 122 nsew signal input
flabel metal2 s 316008 -960 316232 480 0 FreeSans 896 90 0 0 la_data_in[18]
port 123 nsew signal input
flabel metal2 s 321720 -960 321944 480 0 FreeSans 896 90 0 0 la_data_in[19]
port 124 nsew signal input
flabel metal2 s 218904 -960 219128 480 0 FreeSans 896 90 0 0 la_data_in[1]
port 125 nsew signal input
flabel metal2 s 327432 -960 327656 480 0 FreeSans 896 90 0 0 la_data_in[20]
port 126 nsew signal input
flabel metal2 s 333144 -960 333368 480 0 FreeSans 896 90 0 0 la_data_in[21]
port 127 nsew signal input
flabel metal2 s 338856 -960 339080 480 0 FreeSans 896 90 0 0 la_data_in[22]
port 128 nsew signal input
flabel metal2 s 344568 -960 344792 480 0 FreeSans 896 90 0 0 la_data_in[23]
port 129 nsew signal input
flabel metal2 s 350280 -960 350504 480 0 FreeSans 896 90 0 0 la_data_in[24]
port 130 nsew signal input
flabel metal2 s 355992 -960 356216 480 0 FreeSans 896 90 0 0 la_data_in[25]
port 131 nsew signal input
flabel metal2 s 361704 -960 361928 480 0 FreeSans 896 90 0 0 la_data_in[26]
port 132 nsew signal input
flabel metal2 s 367416 -960 367640 480 0 FreeSans 896 90 0 0 la_data_in[27]
port 133 nsew signal input
flabel metal2 s 373128 -960 373352 480 0 FreeSans 896 90 0 0 la_data_in[28]
port 134 nsew signal input
flabel metal2 s 378840 -960 379064 480 0 FreeSans 896 90 0 0 la_data_in[29]
port 135 nsew signal input
flabel metal2 s 224616 -960 224840 480 0 FreeSans 896 90 0 0 la_data_in[2]
port 136 nsew signal input
flabel metal2 s 384552 -960 384776 480 0 FreeSans 896 90 0 0 la_data_in[30]
port 137 nsew signal input
flabel metal2 s 390264 -960 390488 480 0 FreeSans 896 90 0 0 la_data_in[31]
port 138 nsew signal input
flabel metal2 s 395976 -960 396200 480 0 FreeSans 896 90 0 0 la_data_in[32]
port 139 nsew signal input
flabel metal2 s 401688 -960 401912 480 0 FreeSans 896 90 0 0 la_data_in[33]
port 140 nsew signal input
flabel metal2 s 407400 -960 407624 480 0 FreeSans 896 90 0 0 la_data_in[34]
port 141 nsew signal input
flabel metal2 s 413112 -960 413336 480 0 FreeSans 896 90 0 0 la_data_in[35]
port 142 nsew signal input
flabel metal2 s 418824 -960 419048 480 0 FreeSans 896 90 0 0 la_data_in[36]
port 143 nsew signal input
flabel metal2 s 424536 -960 424760 480 0 FreeSans 896 90 0 0 la_data_in[37]
port 144 nsew signal input
flabel metal2 s 430248 -960 430472 480 0 FreeSans 896 90 0 0 la_data_in[38]
port 145 nsew signal input
flabel metal2 s 435960 -960 436184 480 0 FreeSans 896 90 0 0 la_data_in[39]
port 146 nsew signal input
flabel metal2 s 230328 -960 230552 480 0 FreeSans 896 90 0 0 la_data_in[3]
port 147 nsew signal input
flabel metal2 s 441672 -960 441896 480 0 FreeSans 896 90 0 0 la_data_in[40]
port 148 nsew signal input
flabel metal2 s 447384 -960 447608 480 0 FreeSans 896 90 0 0 la_data_in[41]
port 149 nsew signal input
flabel metal2 s 453096 -960 453320 480 0 FreeSans 896 90 0 0 la_data_in[42]
port 150 nsew signal input
flabel metal2 s 458808 -960 459032 480 0 FreeSans 896 90 0 0 la_data_in[43]
port 151 nsew signal input
flabel metal2 s 464520 -960 464744 480 0 FreeSans 896 90 0 0 la_data_in[44]
port 152 nsew signal input
flabel metal2 s 470232 -960 470456 480 0 FreeSans 896 90 0 0 la_data_in[45]
port 153 nsew signal input
flabel metal2 s 475944 -960 476168 480 0 FreeSans 896 90 0 0 la_data_in[46]
port 154 nsew signal input
flabel metal2 s 481656 -960 481880 480 0 FreeSans 896 90 0 0 la_data_in[47]
port 155 nsew signal input
flabel metal2 s 487368 -960 487592 480 0 FreeSans 896 90 0 0 la_data_in[48]
port 156 nsew signal input
flabel metal2 s 493080 -960 493304 480 0 FreeSans 896 90 0 0 la_data_in[49]
port 157 nsew signal input
flabel metal2 s 236040 -960 236264 480 0 FreeSans 896 90 0 0 la_data_in[4]
port 158 nsew signal input
flabel metal2 s 498792 -960 499016 480 0 FreeSans 896 90 0 0 la_data_in[50]
port 159 nsew signal input
flabel metal2 s 504504 -960 504728 480 0 FreeSans 896 90 0 0 la_data_in[51]
port 160 nsew signal input
flabel metal2 s 510216 -960 510440 480 0 FreeSans 896 90 0 0 la_data_in[52]
port 161 nsew signal input
flabel metal2 s 515928 -960 516152 480 0 FreeSans 896 90 0 0 la_data_in[53]
port 162 nsew signal input
flabel metal2 s 521640 -960 521864 480 0 FreeSans 896 90 0 0 la_data_in[54]
port 163 nsew signal input
flabel metal2 s 527352 -960 527576 480 0 FreeSans 896 90 0 0 la_data_in[55]
port 164 nsew signal input
flabel metal2 s 533064 -960 533288 480 0 FreeSans 896 90 0 0 la_data_in[56]
port 165 nsew signal input
flabel metal2 s 538776 -960 539000 480 0 FreeSans 896 90 0 0 la_data_in[57]
port 166 nsew signal input
flabel metal2 s 544488 -960 544712 480 0 FreeSans 896 90 0 0 la_data_in[58]
port 167 nsew signal input
flabel metal2 s 550200 -960 550424 480 0 FreeSans 896 90 0 0 la_data_in[59]
port 168 nsew signal input
flabel metal2 s 241752 -960 241976 480 0 FreeSans 896 90 0 0 la_data_in[5]
port 169 nsew signal input
flabel metal2 s 555912 -960 556136 480 0 FreeSans 896 90 0 0 la_data_in[60]
port 170 nsew signal input
flabel metal2 s 561624 -960 561848 480 0 FreeSans 896 90 0 0 la_data_in[61]
port 171 nsew signal input
flabel metal2 s 567336 -960 567560 480 0 FreeSans 896 90 0 0 la_data_in[62]
port 172 nsew signal input
flabel metal2 s 573048 -960 573272 480 0 FreeSans 896 90 0 0 la_data_in[63]
port 173 nsew signal input
flabel metal2 s 247464 -960 247688 480 0 FreeSans 896 90 0 0 la_data_in[6]
port 174 nsew signal input
flabel metal2 s 253176 -960 253400 480 0 FreeSans 896 90 0 0 la_data_in[7]
port 175 nsew signal input
flabel metal2 s 258888 -960 259112 480 0 FreeSans 896 90 0 0 la_data_in[8]
port 176 nsew signal input
flabel metal2 s 264600 -960 264824 480 0 FreeSans 896 90 0 0 la_data_in[9]
port 177 nsew signal input
flabel metal2 s 215096 -960 215320 480 0 FreeSans 896 90 0 0 la_data_out[0]
port 178 nsew signal tristate
flabel metal2 s 272216 -960 272440 480 0 FreeSans 896 90 0 0 la_data_out[10]
port 179 nsew signal tristate
flabel metal2 s 277928 -960 278152 480 0 FreeSans 896 90 0 0 la_data_out[11]
port 180 nsew signal tristate
flabel metal2 s 283640 -960 283864 480 0 FreeSans 896 90 0 0 la_data_out[12]
port 181 nsew signal tristate
flabel metal2 s 289352 -960 289576 480 0 FreeSans 896 90 0 0 la_data_out[13]
port 182 nsew signal tristate
flabel metal2 s 295064 -960 295288 480 0 FreeSans 896 90 0 0 la_data_out[14]
port 183 nsew signal tristate
flabel metal2 s 300776 -960 301000 480 0 FreeSans 896 90 0 0 la_data_out[15]
port 184 nsew signal tristate
flabel metal2 s 306488 -960 306712 480 0 FreeSans 896 90 0 0 la_data_out[16]
port 185 nsew signal tristate
flabel metal2 s 312200 -960 312424 480 0 FreeSans 896 90 0 0 la_data_out[17]
port 186 nsew signal tristate
flabel metal2 s 317912 -960 318136 480 0 FreeSans 896 90 0 0 la_data_out[18]
port 187 nsew signal tristate
flabel metal2 s 323624 -960 323848 480 0 FreeSans 896 90 0 0 la_data_out[19]
port 188 nsew signal tristate
flabel metal2 s 220808 -960 221032 480 0 FreeSans 896 90 0 0 la_data_out[1]
port 189 nsew signal tristate
flabel metal2 s 329336 -960 329560 480 0 FreeSans 896 90 0 0 la_data_out[20]
port 190 nsew signal tristate
flabel metal2 s 335048 -960 335272 480 0 FreeSans 896 90 0 0 la_data_out[21]
port 191 nsew signal tristate
flabel metal2 s 340760 -960 340984 480 0 FreeSans 896 90 0 0 la_data_out[22]
port 192 nsew signal tristate
flabel metal2 s 346472 -960 346696 480 0 FreeSans 896 90 0 0 la_data_out[23]
port 193 nsew signal tristate
flabel metal2 s 352184 -960 352408 480 0 FreeSans 896 90 0 0 la_data_out[24]
port 194 nsew signal tristate
flabel metal2 s 357896 -960 358120 480 0 FreeSans 896 90 0 0 la_data_out[25]
port 195 nsew signal tristate
flabel metal2 s 363608 -960 363832 480 0 FreeSans 896 90 0 0 la_data_out[26]
port 196 nsew signal tristate
flabel metal2 s 369320 -960 369544 480 0 FreeSans 896 90 0 0 la_data_out[27]
port 197 nsew signal tristate
flabel metal2 s 375032 -960 375256 480 0 FreeSans 896 90 0 0 la_data_out[28]
port 198 nsew signal tristate
flabel metal2 s 380744 -960 380968 480 0 FreeSans 896 90 0 0 la_data_out[29]
port 199 nsew signal tristate
flabel metal2 s 226520 -960 226744 480 0 FreeSans 896 90 0 0 la_data_out[2]
port 200 nsew signal tristate
flabel metal2 s 386456 -960 386680 480 0 FreeSans 896 90 0 0 la_data_out[30]
port 201 nsew signal tristate
flabel metal2 s 392168 -960 392392 480 0 FreeSans 896 90 0 0 la_data_out[31]
port 202 nsew signal tristate
flabel metal2 s 397880 -960 398104 480 0 FreeSans 896 90 0 0 la_data_out[32]
port 203 nsew signal tristate
flabel metal2 s 403592 -960 403816 480 0 FreeSans 896 90 0 0 la_data_out[33]
port 204 nsew signal tristate
flabel metal2 s 409304 -960 409528 480 0 FreeSans 896 90 0 0 la_data_out[34]
port 205 nsew signal tristate
flabel metal2 s 415016 -960 415240 480 0 FreeSans 896 90 0 0 la_data_out[35]
port 206 nsew signal tristate
flabel metal2 s 420728 -960 420952 480 0 FreeSans 896 90 0 0 la_data_out[36]
port 207 nsew signal tristate
flabel metal2 s 426440 -960 426664 480 0 FreeSans 896 90 0 0 la_data_out[37]
port 208 nsew signal tristate
flabel metal2 s 432152 -960 432376 480 0 FreeSans 896 90 0 0 la_data_out[38]
port 209 nsew signal tristate
flabel metal2 s 437864 -960 438088 480 0 FreeSans 896 90 0 0 la_data_out[39]
port 210 nsew signal tristate
flabel metal2 s 232232 -960 232456 480 0 FreeSans 896 90 0 0 la_data_out[3]
port 211 nsew signal tristate
flabel metal2 s 443576 -960 443800 480 0 FreeSans 896 90 0 0 la_data_out[40]
port 212 nsew signal tristate
flabel metal2 s 449288 -960 449512 480 0 FreeSans 896 90 0 0 la_data_out[41]
port 213 nsew signal tristate
flabel metal2 s 455000 -960 455224 480 0 FreeSans 896 90 0 0 la_data_out[42]
port 214 nsew signal tristate
flabel metal2 s 460712 -960 460936 480 0 FreeSans 896 90 0 0 la_data_out[43]
port 215 nsew signal tristate
flabel metal2 s 466424 -960 466648 480 0 FreeSans 896 90 0 0 la_data_out[44]
port 216 nsew signal tristate
flabel metal2 s 472136 -960 472360 480 0 FreeSans 896 90 0 0 la_data_out[45]
port 217 nsew signal tristate
flabel metal2 s 477848 -960 478072 480 0 FreeSans 896 90 0 0 la_data_out[46]
port 218 nsew signal tristate
flabel metal2 s 483560 -960 483784 480 0 FreeSans 896 90 0 0 la_data_out[47]
port 219 nsew signal tristate
flabel metal2 s 489272 -960 489496 480 0 FreeSans 896 90 0 0 la_data_out[48]
port 220 nsew signal tristate
flabel metal2 s 494984 -960 495208 480 0 FreeSans 896 90 0 0 la_data_out[49]
port 221 nsew signal tristate
flabel metal2 s 237944 -960 238168 480 0 FreeSans 896 90 0 0 la_data_out[4]
port 222 nsew signal tristate
flabel metal2 s 500696 -960 500920 480 0 FreeSans 896 90 0 0 la_data_out[50]
port 223 nsew signal tristate
flabel metal2 s 506408 -960 506632 480 0 FreeSans 896 90 0 0 la_data_out[51]
port 224 nsew signal tristate
flabel metal2 s 512120 -960 512344 480 0 FreeSans 896 90 0 0 la_data_out[52]
port 225 nsew signal tristate
flabel metal2 s 517832 -960 518056 480 0 FreeSans 896 90 0 0 la_data_out[53]
port 226 nsew signal tristate
flabel metal2 s 523544 -960 523768 480 0 FreeSans 896 90 0 0 la_data_out[54]
port 227 nsew signal tristate
flabel metal2 s 529256 -960 529480 480 0 FreeSans 896 90 0 0 la_data_out[55]
port 228 nsew signal tristate
flabel metal2 s 534968 -960 535192 480 0 FreeSans 896 90 0 0 la_data_out[56]
port 229 nsew signal tristate
flabel metal2 s 540680 -960 540904 480 0 FreeSans 896 90 0 0 la_data_out[57]
port 230 nsew signal tristate
flabel metal2 s 546392 -960 546616 480 0 FreeSans 896 90 0 0 la_data_out[58]
port 231 nsew signal tristate
flabel metal2 s 552104 -960 552328 480 0 FreeSans 896 90 0 0 la_data_out[59]
port 232 nsew signal tristate
flabel metal2 s 243656 -960 243880 480 0 FreeSans 896 90 0 0 la_data_out[5]
port 233 nsew signal tristate
flabel metal2 s 557816 -960 558040 480 0 FreeSans 896 90 0 0 la_data_out[60]
port 234 nsew signal tristate
flabel metal2 s 563528 -960 563752 480 0 FreeSans 896 90 0 0 la_data_out[61]
port 235 nsew signal tristate
flabel metal2 s 569240 -960 569464 480 0 FreeSans 896 90 0 0 la_data_out[62]
port 236 nsew signal tristate
flabel metal2 s 574952 -960 575176 480 0 FreeSans 896 90 0 0 la_data_out[63]
port 237 nsew signal tristate
flabel metal2 s 249368 -960 249592 480 0 FreeSans 896 90 0 0 la_data_out[6]
port 238 nsew signal tristate
flabel metal2 s 255080 -960 255304 480 0 FreeSans 896 90 0 0 la_data_out[7]
port 239 nsew signal tristate
flabel metal2 s 260792 -960 261016 480 0 FreeSans 896 90 0 0 la_data_out[8]
port 240 nsew signal tristate
flabel metal2 s 266504 -960 266728 480 0 FreeSans 896 90 0 0 la_data_out[9]
port 241 nsew signal tristate
flabel metal2 s 217000 -960 217224 480 0 FreeSans 896 90 0 0 la_oenb[0]
port 242 nsew signal input
flabel metal2 s 274120 -960 274344 480 0 FreeSans 896 90 0 0 la_oenb[10]
port 243 nsew signal input
flabel metal2 s 279832 -960 280056 480 0 FreeSans 896 90 0 0 la_oenb[11]
port 244 nsew signal input
flabel metal2 s 285544 -960 285768 480 0 FreeSans 896 90 0 0 la_oenb[12]
port 245 nsew signal input
flabel metal2 s 291256 -960 291480 480 0 FreeSans 896 90 0 0 la_oenb[13]
port 246 nsew signal input
flabel metal2 s 296968 -960 297192 480 0 FreeSans 896 90 0 0 la_oenb[14]
port 247 nsew signal input
flabel metal2 s 302680 -960 302904 480 0 FreeSans 896 90 0 0 la_oenb[15]
port 248 nsew signal input
flabel metal2 s 308392 -960 308616 480 0 FreeSans 896 90 0 0 la_oenb[16]
port 249 nsew signal input
flabel metal2 s 314104 -960 314328 480 0 FreeSans 896 90 0 0 la_oenb[17]
port 250 nsew signal input
flabel metal2 s 319816 -960 320040 480 0 FreeSans 896 90 0 0 la_oenb[18]
port 251 nsew signal input
flabel metal2 s 325528 -960 325752 480 0 FreeSans 896 90 0 0 la_oenb[19]
port 252 nsew signal input
flabel metal2 s 222712 -960 222936 480 0 FreeSans 896 90 0 0 la_oenb[1]
port 253 nsew signal input
flabel metal2 s 331240 -960 331464 480 0 FreeSans 896 90 0 0 la_oenb[20]
port 254 nsew signal input
flabel metal2 s 336952 -960 337176 480 0 FreeSans 896 90 0 0 la_oenb[21]
port 255 nsew signal input
flabel metal2 s 342664 -960 342888 480 0 FreeSans 896 90 0 0 la_oenb[22]
port 256 nsew signal input
flabel metal2 s 348376 -960 348600 480 0 FreeSans 896 90 0 0 la_oenb[23]
port 257 nsew signal input
flabel metal2 s 354088 -960 354312 480 0 FreeSans 896 90 0 0 la_oenb[24]
port 258 nsew signal input
flabel metal2 s 359800 -960 360024 480 0 FreeSans 896 90 0 0 la_oenb[25]
port 259 nsew signal input
flabel metal2 s 365512 -960 365736 480 0 FreeSans 896 90 0 0 la_oenb[26]
port 260 nsew signal input
flabel metal2 s 371224 -960 371448 480 0 FreeSans 896 90 0 0 la_oenb[27]
port 261 nsew signal input
flabel metal2 s 376936 -960 377160 480 0 FreeSans 896 90 0 0 la_oenb[28]
port 262 nsew signal input
flabel metal2 s 382648 -960 382872 480 0 FreeSans 896 90 0 0 la_oenb[29]
port 263 nsew signal input
flabel metal2 s 228424 -960 228648 480 0 FreeSans 896 90 0 0 la_oenb[2]
port 264 nsew signal input
flabel metal2 s 388360 -960 388584 480 0 FreeSans 896 90 0 0 la_oenb[30]
port 265 nsew signal input
flabel metal2 s 394072 -960 394296 480 0 FreeSans 896 90 0 0 la_oenb[31]
port 266 nsew signal input
flabel metal2 s 399784 -960 400008 480 0 FreeSans 896 90 0 0 la_oenb[32]
port 267 nsew signal input
flabel metal2 s 405496 -960 405720 480 0 FreeSans 896 90 0 0 la_oenb[33]
port 268 nsew signal input
flabel metal2 s 411208 -960 411432 480 0 FreeSans 896 90 0 0 la_oenb[34]
port 269 nsew signal input
flabel metal2 s 416920 -960 417144 480 0 FreeSans 896 90 0 0 la_oenb[35]
port 270 nsew signal input
flabel metal2 s 422632 -960 422856 480 0 FreeSans 896 90 0 0 la_oenb[36]
port 271 nsew signal input
flabel metal2 s 428344 -960 428568 480 0 FreeSans 896 90 0 0 la_oenb[37]
port 272 nsew signal input
flabel metal2 s 434056 -960 434280 480 0 FreeSans 896 90 0 0 la_oenb[38]
port 273 nsew signal input
flabel metal2 s 439768 -960 439992 480 0 FreeSans 896 90 0 0 la_oenb[39]
port 274 nsew signal input
flabel metal2 s 234136 -960 234360 480 0 FreeSans 896 90 0 0 la_oenb[3]
port 275 nsew signal input
flabel metal2 s 445480 -960 445704 480 0 FreeSans 896 90 0 0 la_oenb[40]
port 276 nsew signal input
flabel metal2 s 451192 -960 451416 480 0 FreeSans 896 90 0 0 la_oenb[41]
port 277 nsew signal input
flabel metal2 s 456904 -960 457128 480 0 FreeSans 896 90 0 0 la_oenb[42]
port 278 nsew signal input
flabel metal2 s 462616 -960 462840 480 0 FreeSans 896 90 0 0 la_oenb[43]
port 279 nsew signal input
flabel metal2 s 468328 -960 468552 480 0 FreeSans 896 90 0 0 la_oenb[44]
port 280 nsew signal input
flabel metal2 s 474040 -960 474264 480 0 FreeSans 896 90 0 0 la_oenb[45]
port 281 nsew signal input
flabel metal2 s 479752 -960 479976 480 0 FreeSans 896 90 0 0 la_oenb[46]
port 282 nsew signal input
flabel metal2 s 485464 -960 485688 480 0 FreeSans 896 90 0 0 la_oenb[47]
port 283 nsew signal input
flabel metal2 s 491176 -960 491400 480 0 FreeSans 896 90 0 0 la_oenb[48]
port 284 nsew signal input
flabel metal2 s 496888 -960 497112 480 0 FreeSans 896 90 0 0 la_oenb[49]
port 285 nsew signal input
flabel metal2 s 239848 -960 240072 480 0 FreeSans 896 90 0 0 la_oenb[4]
port 286 nsew signal input
flabel metal2 s 502600 -960 502824 480 0 FreeSans 896 90 0 0 la_oenb[50]
port 287 nsew signal input
flabel metal2 s 508312 -960 508536 480 0 FreeSans 896 90 0 0 la_oenb[51]
port 288 nsew signal input
flabel metal2 s 514024 -960 514248 480 0 FreeSans 896 90 0 0 la_oenb[52]
port 289 nsew signal input
flabel metal2 s 519736 -960 519960 480 0 FreeSans 896 90 0 0 la_oenb[53]
port 290 nsew signal input
flabel metal2 s 525448 -960 525672 480 0 FreeSans 896 90 0 0 la_oenb[54]
port 291 nsew signal input
flabel metal2 s 531160 -960 531384 480 0 FreeSans 896 90 0 0 la_oenb[55]
port 292 nsew signal input
flabel metal2 s 536872 -960 537096 480 0 FreeSans 896 90 0 0 la_oenb[56]
port 293 nsew signal input
flabel metal2 s 542584 -960 542808 480 0 FreeSans 896 90 0 0 la_oenb[57]
port 294 nsew signal input
flabel metal2 s 548296 -960 548520 480 0 FreeSans 896 90 0 0 la_oenb[58]
port 295 nsew signal input
flabel metal2 s 554008 -960 554232 480 0 FreeSans 896 90 0 0 la_oenb[59]
port 296 nsew signal input
flabel metal2 s 245560 -960 245784 480 0 FreeSans 896 90 0 0 la_oenb[5]
port 297 nsew signal input
flabel metal2 s 559720 -960 559944 480 0 FreeSans 896 90 0 0 la_oenb[60]
port 298 nsew signal input
flabel metal2 s 565432 -960 565656 480 0 FreeSans 896 90 0 0 la_oenb[61]
port 299 nsew signal input
flabel metal2 s 571144 -960 571368 480 0 FreeSans 896 90 0 0 la_oenb[62]
port 300 nsew signal input
flabel metal2 s 576856 -960 577080 480 0 FreeSans 896 90 0 0 la_oenb[63]
port 301 nsew signal input
flabel metal2 s 251272 -960 251496 480 0 FreeSans 896 90 0 0 la_oenb[6]
port 302 nsew signal input
flabel metal2 s 256984 -960 257208 480 0 FreeSans 896 90 0 0 la_oenb[7]
port 303 nsew signal input
flabel metal2 s 262696 -960 262920 480 0 FreeSans 896 90 0 0 la_oenb[8]
port 304 nsew signal input
flabel metal2 s 268408 -960 268632 480 0 FreeSans 896 90 0 0 la_oenb[9]
port 305 nsew signal input
flabel metal2 s 578760 -960 578984 480 0 FreeSans 896 90 0 0 user_clock2
port 306 nsew signal input
flabel metal2 s 580664 -960 580888 480 0 FreeSans 896 90 0 0 user_irq[0]
port 307 nsew signal tristate
flabel metal2 s 582568 -960 582792 480 0 FreeSans 896 90 0 0 user_irq[1]
port 308 nsew signal tristate
flabel metal2 s 584472 -960 584696 480 0 FreeSans 896 90 0 0 user_irq[2]
port 309 nsew signal tristate
flabel metal4 s -956 -684 -336 597308 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -956 -684 597020 -64 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -956 596688 597020 597308 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 596400 -684 597020 597308 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 3154 -1644 3774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 21154 -1644 21774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 39154 -1644 39774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 57154 -1644 57774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 75154 -1644 75774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 93154 -1644 93774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 111154 -1644 111774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 129154 -1644 129774 32890 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 129154 527750 129774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 147154 -1644 147774 32890 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 147154 527750 147774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 165154 -1644 165774 32890 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 165154 527750 165774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 183154 -1644 183774 32890 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 183154 527750 183774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 201154 -1644 201774 32890 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 201154 527750 201774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 219154 -1644 219774 32890 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 219154 527750 219774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 237154 -1644 237774 32890 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 237154 527750 237774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 255154 -1644 255774 32890 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 255154 527750 255774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 273154 -1644 273774 32890 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 273154 527750 273774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 291154 -1644 291774 32890 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 291154 527750 291774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 309154 -1644 309774 32890 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 309154 527750 309774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 327154 -1644 327774 32890 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 327154 527750 327774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 345154 -1644 345774 32890 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 345154 527750 345774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 363154 -1644 363774 32890 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 363154 527750 363774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 381154 -1644 381774 32890 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 381154 527750 381774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 399154 -1644 399774 32890 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 399154 527750 399774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 417154 -1644 417774 32890 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 417154 527750 417774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 435154 -1644 435774 32890 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 435154 527750 435774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 453154 -1644 453774 31020 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 453154 528388 453774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 471154 -1644 471774 32890 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 471154 527750 471774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 489154 -1644 489774 32890 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 489154 527750 489774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 507154 -1644 507774 32890 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 507154 527750 507774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 525154 -1644 525774 32890 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 525154 527750 525774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 543154 -1644 543774 32890 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 543154 527750 543774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 561154 -1644 561774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 579154 -1644 579774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 3826 597980 4446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 21826 597980 22446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 39826 597980 40446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 57826 597980 58446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 75826 597980 76446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 93826 597980 94446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 111826 597980 112446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 129826 597980 130446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 147826 597980 148446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 165826 597980 166446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 183826 597980 184446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 201826 597980 202446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 219826 597980 220446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 237826 597980 238446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 255826 597980 256446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 273826 597980 274446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 291826 597980 292446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 309826 597980 310446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 327826 597980 328446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 345826 597980 346446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 363826 597980 364446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 381826 597980 382446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 399826 597980 400446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 417826 597980 418446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 435826 597980 436446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 453826 597980 454446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 471826 597980 472446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 489826 597980 490446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 507826 597980 508446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 525826 597980 526446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 543826 597980 544446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 561826 597980 562446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 579826 597980 580446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s -1916 -1644 -1296 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 -1644 597980 -1024 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 597648 597980 598268 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 597360 -1644 597980 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 6874 -1644 7494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 24874 -1644 25494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 42874 -1644 43494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 60874 -1644 61494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 78874 -1644 79494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 96874 -1644 97494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 114874 -1644 115494 32890 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 114874 527750 115494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 132874 -1644 133494 32890 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 132874 527750 133494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 150874 -1644 151494 32890 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 150874 527750 151494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 168874 -1644 169494 32890 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 168874 527750 169494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 186874 -1644 187494 32890 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 186874 527750 187494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 204874 -1644 205494 32890 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 204874 527750 205494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 222874 -1644 223494 31020 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 222874 528388 223494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 240874 -1644 241494 32890 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 240874 527750 241494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 258874 -1644 259494 32890 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 258874 527750 259494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 276874 -1644 277494 32890 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 276874 527750 277494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 294874 -1644 295494 32890 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 294874 527750 295494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 312874 -1644 313494 32890 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 312874 527750 313494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 330874 -1644 331494 31020 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 330874 528388 331494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 348874 -1644 349494 32890 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 348874 527750 349494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 366874 -1644 367494 32890 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 366874 527750 367494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 384874 -1644 385494 32890 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 384874 527750 385494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 402874 -1644 403494 32890 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 402874 527750 403494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 420874 -1644 421494 32890 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 420874 527750 421494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 438874 -1644 439494 32890 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 438874 527750 439494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 456874 -1644 457494 32890 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 456874 527750 457494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 474874 -1644 475494 32890 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 474874 527750 475494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 492874 -1644 493494 32890 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 492874 527750 493494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 510874 -1644 511494 32890 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 510874 527750 511494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 528874 -1644 529494 32890 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 528874 527750 529494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 546874 -1644 547494 32890 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 546874 527750 547494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 564874 -1644 565494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 582874 -1644 583494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 9826 597980 10446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 27826 597980 28446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 45826 597980 46446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 63826 597980 64446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 81826 597980 82446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 99826 597980 100446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 117826 597980 118446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 135826 597980 136446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 153826 597980 154446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 171826 597980 172446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 189826 597980 190446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 207826 597980 208446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 225826 597980 226446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 243826 597980 244446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 261826 597980 262446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 279826 597980 280446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 297826 597980 298446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 315826 597980 316446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 333826 597980 334446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 351826 597980 352446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 369826 597980 370446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 387826 597980 388446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 405826 597980 406446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 423826 597980 424446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 441826 597980 442446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 459826 597980 460446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 477826 597980 478446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 495826 597980 496446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 513826 597980 514446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 531826 597980 532446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 549826 597980 550446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 567826 597980 568446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 585826 597980 586446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal2 s 11368 -960 11592 480 0 FreeSans 896 90 0 0 wb_clk_i
port 312 nsew signal input
flabel metal2 s 13272 -960 13496 480 0 FreeSans 896 90 0 0 wb_rst_i
port 313 nsew signal input
flabel metal2 s 15176 -960 15400 480 0 FreeSans 896 90 0 0 wbs_ack_o
port 314 nsew signal tristate
flabel metal2 s 22792 -960 23016 480 0 FreeSans 896 90 0 0 wbs_adr_i[0]
port 315 nsew signal input
flabel metal2 s 87528 -960 87752 480 0 FreeSans 896 90 0 0 wbs_adr_i[10]
port 316 nsew signal input
flabel metal2 s 93240 -960 93464 480 0 FreeSans 896 90 0 0 wbs_adr_i[11]
port 317 nsew signal input
flabel metal2 s 98952 -960 99176 480 0 FreeSans 896 90 0 0 wbs_adr_i[12]
port 318 nsew signal input
flabel metal2 s 104664 -960 104888 480 0 FreeSans 896 90 0 0 wbs_adr_i[13]
port 319 nsew signal input
flabel metal2 s 110376 -960 110600 480 0 FreeSans 896 90 0 0 wbs_adr_i[14]
port 320 nsew signal input
flabel metal2 s 116088 -960 116312 480 0 FreeSans 896 90 0 0 wbs_adr_i[15]
port 321 nsew signal input
flabel metal2 s 121800 -960 122024 480 0 FreeSans 896 90 0 0 wbs_adr_i[16]
port 322 nsew signal input
flabel metal2 s 127512 -960 127736 480 0 FreeSans 896 90 0 0 wbs_adr_i[17]
port 323 nsew signal input
flabel metal2 s 133224 -960 133448 480 0 FreeSans 896 90 0 0 wbs_adr_i[18]
port 324 nsew signal input
flabel metal2 s 138936 -960 139160 480 0 FreeSans 896 90 0 0 wbs_adr_i[19]
port 325 nsew signal input
flabel metal2 s 30408 -960 30632 480 0 FreeSans 896 90 0 0 wbs_adr_i[1]
port 326 nsew signal input
flabel metal2 s 144648 -960 144872 480 0 FreeSans 896 90 0 0 wbs_adr_i[20]
port 327 nsew signal input
flabel metal2 s 150360 -960 150584 480 0 FreeSans 896 90 0 0 wbs_adr_i[21]
port 328 nsew signal input
flabel metal2 s 156072 -960 156296 480 0 FreeSans 896 90 0 0 wbs_adr_i[22]
port 329 nsew signal input
flabel metal2 s 161784 -960 162008 480 0 FreeSans 896 90 0 0 wbs_adr_i[23]
port 330 nsew signal input
flabel metal2 s 167496 -960 167720 480 0 FreeSans 896 90 0 0 wbs_adr_i[24]
port 331 nsew signal input
flabel metal2 s 173208 -960 173432 480 0 FreeSans 896 90 0 0 wbs_adr_i[25]
port 332 nsew signal input
flabel metal2 s 178920 -960 179144 480 0 FreeSans 896 90 0 0 wbs_adr_i[26]
port 333 nsew signal input
flabel metal2 s 184632 -960 184856 480 0 FreeSans 896 90 0 0 wbs_adr_i[27]
port 334 nsew signal input
flabel metal2 s 190344 -960 190568 480 0 FreeSans 896 90 0 0 wbs_adr_i[28]
port 335 nsew signal input
flabel metal2 s 196056 -960 196280 480 0 FreeSans 896 90 0 0 wbs_adr_i[29]
port 336 nsew signal input
flabel metal2 s 38024 -960 38248 480 0 FreeSans 896 90 0 0 wbs_adr_i[2]
port 337 nsew signal input
flabel metal2 s 201768 -960 201992 480 0 FreeSans 896 90 0 0 wbs_adr_i[30]
port 338 nsew signal input
flabel metal2 s 207480 -960 207704 480 0 FreeSans 896 90 0 0 wbs_adr_i[31]
port 339 nsew signal input
flabel metal2 s 45640 -960 45864 480 0 FreeSans 896 90 0 0 wbs_adr_i[3]
port 340 nsew signal input
flabel metal2 s 53256 -960 53480 480 0 FreeSans 896 90 0 0 wbs_adr_i[4]
port 341 nsew signal input
flabel metal2 s 58968 -960 59192 480 0 FreeSans 896 90 0 0 wbs_adr_i[5]
port 342 nsew signal input
flabel metal2 s 64680 -960 64904 480 0 FreeSans 896 90 0 0 wbs_adr_i[6]
port 343 nsew signal input
flabel metal2 s 70392 -960 70616 480 0 FreeSans 896 90 0 0 wbs_adr_i[7]
port 344 nsew signal input
flabel metal2 s 76104 -960 76328 480 0 FreeSans 896 90 0 0 wbs_adr_i[8]
port 345 nsew signal input
flabel metal2 s 81816 -960 82040 480 0 FreeSans 896 90 0 0 wbs_adr_i[9]
port 346 nsew signal input
flabel metal2 s 17080 -960 17304 480 0 FreeSans 896 90 0 0 wbs_cyc_i
port 347 nsew signal input
flabel metal2 s 24696 -960 24920 480 0 FreeSans 896 90 0 0 wbs_dat_i[0]
port 348 nsew signal input
flabel metal2 s 89432 -960 89656 480 0 FreeSans 896 90 0 0 wbs_dat_i[10]
port 349 nsew signal input
flabel metal2 s 95144 -960 95368 480 0 FreeSans 896 90 0 0 wbs_dat_i[11]
port 350 nsew signal input
flabel metal2 s 100856 -960 101080 480 0 FreeSans 896 90 0 0 wbs_dat_i[12]
port 351 nsew signal input
flabel metal2 s 106568 -960 106792 480 0 FreeSans 896 90 0 0 wbs_dat_i[13]
port 352 nsew signal input
flabel metal2 s 112280 -960 112504 480 0 FreeSans 896 90 0 0 wbs_dat_i[14]
port 353 nsew signal input
flabel metal2 s 117992 -960 118216 480 0 FreeSans 896 90 0 0 wbs_dat_i[15]
port 354 nsew signal input
flabel metal2 s 123704 -960 123928 480 0 FreeSans 896 90 0 0 wbs_dat_i[16]
port 355 nsew signal input
flabel metal2 s 129416 -960 129640 480 0 FreeSans 896 90 0 0 wbs_dat_i[17]
port 356 nsew signal input
flabel metal2 s 135128 -960 135352 480 0 FreeSans 896 90 0 0 wbs_dat_i[18]
port 357 nsew signal input
flabel metal2 s 140840 -960 141064 480 0 FreeSans 896 90 0 0 wbs_dat_i[19]
port 358 nsew signal input
flabel metal2 s 32312 -960 32536 480 0 FreeSans 896 90 0 0 wbs_dat_i[1]
port 359 nsew signal input
flabel metal2 s 146552 -960 146776 480 0 FreeSans 896 90 0 0 wbs_dat_i[20]
port 360 nsew signal input
flabel metal2 s 152264 -960 152488 480 0 FreeSans 896 90 0 0 wbs_dat_i[21]
port 361 nsew signal input
flabel metal2 s 157976 -960 158200 480 0 FreeSans 896 90 0 0 wbs_dat_i[22]
port 362 nsew signal input
flabel metal2 s 163688 -960 163912 480 0 FreeSans 896 90 0 0 wbs_dat_i[23]
port 363 nsew signal input
flabel metal2 s 169400 -960 169624 480 0 FreeSans 896 90 0 0 wbs_dat_i[24]
port 364 nsew signal input
flabel metal2 s 175112 -960 175336 480 0 FreeSans 896 90 0 0 wbs_dat_i[25]
port 365 nsew signal input
flabel metal2 s 180824 -960 181048 480 0 FreeSans 896 90 0 0 wbs_dat_i[26]
port 366 nsew signal input
flabel metal2 s 186536 -960 186760 480 0 FreeSans 896 90 0 0 wbs_dat_i[27]
port 367 nsew signal input
flabel metal2 s 192248 -960 192472 480 0 FreeSans 896 90 0 0 wbs_dat_i[28]
port 368 nsew signal input
flabel metal2 s 197960 -960 198184 480 0 FreeSans 896 90 0 0 wbs_dat_i[29]
port 369 nsew signal input
flabel metal2 s 39928 -960 40152 480 0 FreeSans 896 90 0 0 wbs_dat_i[2]
port 370 nsew signal input
flabel metal2 s 203672 -960 203896 480 0 FreeSans 896 90 0 0 wbs_dat_i[30]
port 371 nsew signal input
flabel metal2 s 209384 -960 209608 480 0 FreeSans 896 90 0 0 wbs_dat_i[31]
port 372 nsew signal input
flabel metal2 s 47544 -960 47768 480 0 FreeSans 896 90 0 0 wbs_dat_i[3]
port 373 nsew signal input
flabel metal2 s 55160 -960 55384 480 0 FreeSans 896 90 0 0 wbs_dat_i[4]
port 374 nsew signal input
flabel metal2 s 60872 -960 61096 480 0 FreeSans 896 90 0 0 wbs_dat_i[5]
port 375 nsew signal input
flabel metal2 s 66584 -960 66808 480 0 FreeSans 896 90 0 0 wbs_dat_i[6]
port 376 nsew signal input
flabel metal2 s 72296 -960 72520 480 0 FreeSans 896 90 0 0 wbs_dat_i[7]
port 377 nsew signal input
flabel metal2 s 78008 -960 78232 480 0 FreeSans 896 90 0 0 wbs_dat_i[8]
port 378 nsew signal input
flabel metal2 s 83720 -960 83944 480 0 FreeSans 896 90 0 0 wbs_dat_i[9]
port 379 nsew signal input
flabel metal2 s 26600 -960 26824 480 0 FreeSans 896 90 0 0 wbs_dat_o[0]
port 380 nsew signal tristate
flabel metal2 s 91336 -960 91560 480 0 FreeSans 896 90 0 0 wbs_dat_o[10]
port 381 nsew signal tristate
flabel metal2 s 97048 -960 97272 480 0 FreeSans 896 90 0 0 wbs_dat_o[11]
port 382 nsew signal tristate
flabel metal2 s 102760 -960 102984 480 0 FreeSans 896 90 0 0 wbs_dat_o[12]
port 383 nsew signal tristate
flabel metal2 s 108472 -960 108696 480 0 FreeSans 896 90 0 0 wbs_dat_o[13]
port 384 nsew signal tristate
flabel metal2 s 114184 -960 114408 480 0 FreeSans 896 90 0 0 wbs_dat_o[14]
port 385 nsew signal tristate
flabel metal2 s 119896 -960 120120 480 0 FreeSans 896 90 0 0 wbs_dat_o[15]
port 386 nsew signal tristate
flabel metal2 s 125608 -960 125832 480 0 FreeSans 896 90 0 0 wbs_dat_o[16]
port 387 nsew signal tristate
flabel metal2 s 131320 -960 131544 480 0 FreeSans 896 90 0 0 wbs_dat_o[17]
port 388 nsew signal tristate
flabel metal2 s 137032 -960 137256 480 0 FreeSans 896 90 0 0 wbs_dat_o[18]
port 389 nsew signal tristate
flabel metal2 s 142744 -960 142968 480 0 FreeSans 896 90 0 0 wbs_dat_o[19]
port 390 nsew signal tristate
flabel metal2 s 34216 -960 34440 480 0 FreeSans 896 90 0 0 wbs_dat_o[1]
port 391 nsew signal tristate
flabel metal2 s 148456 -960 148680 480 0 FreeSans 896 90 0 0 wbs_dat_o[20]
port 392 nsew signal tristate
flabel metal2 s 154168 -960 154392 480 0 FreeSans 896 90 0 0 wbs_dat_o[21]
port 393 nsew signal tristate
flabel metal2 s 159880 -960 160104 480 0 FreeSans 896 90 0 0 wbs_dat_o[22]
port 394 nsew signal tristate
flabel metal2 s 165592 -960 165816 480 0 FreeSans 896 90 0 0 wbs_dat_o[23]
port 395 nsew signal tristate
flabel metal2 s 171304 -960 171528 480 0 FreeSans 896 90 0 0 wbs_dat_o[24]
port 396 nsew signal tristate
flabel metal2 s 177016 -960 177240 480 0 FreeSans 896 90 0 0 wbs_dat_o[25]
port 397 nsew signal tristate
flabel metal2 s 182728 -960 182952 480 0 FreeSans 896 90 0 0 wbs_dat_o[26]
port 398 nsew signal tristate
flabel metal2 s 188440 -960 188664 480 0 FreeSans 896 90 0 0 wbs_dat_o[27]
port 399 nsew signal tristate
flabel metal2 s 194152 -960 194376 480 0 FreeSans 896 90 0 0 wbs_dat_o[28]
port 400 nsew signal tristate
flabel metal2 s 199864 -960 200088 480 0 FreeSans 896 90 0 0 wbs_dat_o[29]
port 401 nsew signal tristate
flabel metal2 s 41832 -960 42056 480 0 FreeSans 896 90 0 0 wbs_dat_o[2]
port 402 nsew signal tristate
flabel metal2 s 205576 -960 205800 480 0 FreeSans 896 90 0 0 wbs_dat_o[30]
port 403 nsew signal tristate
flabel metal2 s 211288 -960 211512 480 0 FreeSans 896 90 0 0 wbs_dat_o[31]
port 404 nsew signal tristate
flabel metal2 s 49448 -960 49672 480 0 FreeSans 896 90 0 0 wbs_dat_o[3]
port 405 nsew signal tristate
flabel metal2 s 57064 -960 57288 480 0 FreeSans 896 90 0 0 wbs_dat_o[4]
port 406 nsew signal tristate
flabel metal2 s 62776 -960 63000 480 0 FreeSans 896 90 0 0 wbs_dat_o[5]
port 407 nsew signal tristate
flabel metal2 s 68488 -960 68712 480 0 FreeSans 896 90 0 0 wbs_dat_o[6]
port 408 nsew signal tristate
flabel metal2 s 74200 -960 74424 480 0 FreeSans 896 90 0 0 wbs_dat_o[7]
port 409 nsew signal tristate
flabel metal2 s 79912 -960 80136 480 0 FreeSans 896 90 0 0 wbs_dat_o[8]
port 410 nsew signal tristate
flabel metal2 s 85624 -960 85848 480 0 FreeSans 896 90 0 0 wbs_dat_o[9]
port 411 nsew signal tristate
flabel metal2 s 28504 -960 28728 480 0 FreeSans 896 90 0 0 wbs_sel_i[0]
port 412 nsew signal input
flabel metal2 s 36120 -960 36344 480 0 FreeSans 896 90 0 0 wbs_sel_i[1]
port 413 nsew signal input
flabel metal2 s 43736 -960 43960 480 0 FreeSans 896 90 0 0 wbs_sel_i[2]
port 414 nsew signal input
flabel metal2 s 51352 -960 51576 480 0 FreeSans 896 90 0 0 wbs_sel_i[3]
port 415 nsew signal input
flabel metal2 s 18984 -960 19208 480 0 FreeSans 896 90 0 0 wbs_stb_i
port 416 nsew signal input
flabel metal2 s 20888 -960 21112 480 0 FreeSans 896 90 0 0 wbs_we_i
port 417 nsew signal input
rlabel via4 546190 526265 546190 526265 0 vdd
rlabel via4 530830 514322 530830 514322 0 vss
rlabel metal2 11592 2310 11592 2310 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 596040 596040
<< end >>
