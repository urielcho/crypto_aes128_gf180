magic
tech gf180mcuC
magscale 1 5
timestamp 1670226993
<< obsm1 >>
rect 672 1471 249312 248345
<< metal2 >>
rect 1680 249600 1736 249900
rect 4368 249600 4424 249900
rect 7056 249600 7112 249900
rect 9408 249600 9464 249900
rect 12096 249600 12152 249900
rect 14784 249600 14840 249900
rect 17472 249600 17528 249900
rect 19824 249600 19880 249900
rect 22512 249600 22568 249900
rect 25200 249600 25256 249900
rect 27888 249600 27944 249900
rect 30240 249600 30296 249900
rect 32928 249600 32984 249900
rect 35616 249600 35672 249900
rect 38304 249600 38360 249900
rect 40656 249600 40712 249900
rect 43344 249600 43400 249900
rect 46032 249600 46088 249900
rect 48384 249600 48440 249900
rect 51072 249600 51128 249900
rect 53760 249600 53816 249900
rect 56448 249600 56504 249900
rect 58800 249600 58856 249900
rect 61488 249600 61544 249900
rect 64176 249600 64232 249900
rect 66864 249600 66920 249900
rect 69216 249600 69272 249900
rect 71904 249600 71960 249900
rect 74592 249600 74648 249900
rect 76944 249600 77000 249900
rect 79632 249600 79688 249900
rect 82320 249600 82376 249900
rect 85008 249600 85064 249900
rect 87360 249600 87416 249900
rect 90048 249600 90104 249900
rect 92736 249600 92792 249900
rect 95424 249600 95480 249900
rect 97776 249600 97832 249900
rect 100464 249600 100520 249900
rect 103152 249600 103208 249900
rect 105504 249600 105560 249900
rect 108192 249600 108248 249900
rect 110880 249600 110936 249900
rect 113568 249600 113624 249900
rect 115920 249600 115976 249900
rect 118608 249600 118664 249900
rect 121296 249600 121352 249900
rect 123984 249600 124040 249900
rect 126336 249600 126392 249900
rect 129024 249600 129080 249900
rect 131712 249600 131768 249900
rect 134400 249600 134456 249900
rect 136752 249600 136808 249900
rect 139440 249600 139496 249900
rect 142128 249600 142184 249900
rect 144480 249600 144536 249900
rect 147168 249600 147224 249900
rect 149856 249600 149912 249900
rect 152544 249600 152600 249900
rect 154896 249600 154952 249900
rect 157584 249600 157640 249900
rect 160272 249600 160328 249900
rect 162960 249600 163016 249900
rect 165312 249600 165368 249900
rect 168000 249600 168056 249900
rect 170688 249600 170744 249900
rect 173040 249600 173096 249900
rect 175728 249600 175784 249900
rect 178416 249600 178472 249900
rect 181104 249600 181160 249900
rect 183456 249600 183512 249900
rect 186144 249600 186200 249900
rect 188832 249600 188888 249900
rect 191520 249600 191576 249900
rect 193872 249600 193928 249900
rect 196560 249600 196616 249900
rect 199248 249600 199304 249900
rect 201600 249600 201656 249900
rect 204288 249600 204344 249900
rect 206976 249600 207032 249900
rect 209664 249600 209720 249900
rect 212016 249600 212072 249900
rect 214704 249600 214760 249900
rect 217392 249600 217448 249900
rect 220080 249600 220136 249900
rect 222432 249600 222488 249900
rect 225120 249600 225176 249900
rect 227808 249600 227864 249900
rect 230496 249600 230552 249900
rect 232848 249600 232904 249900
rect 235536 249600 235592 249900
rect 238224 249600 238280 249900
rect 240576 249600 240632 249900
rect 243264 249600 243320 249900
rect 245952 249600 246008 249900
rect 248640 249600 248696 249900
rect 0 100 56 400
rect 2352 100 2408 400
rect 5040 100 5096 400
rect 7728 100 7784 400
rect 10080 100 10136 400
rect 12768 100 12824 400
rect 15456 100 15512 400
rect 18144 100 18200 400
rect 20496 100 20552 400
rect 23184 100 23240 400
rect 25872 100 25928 400
rect 28560 100 28616 400
rect 30912 100 30968 400
rect 33600 100 33656 400
rect 36288 100 36344 400
rect 38640 100 38696 400
rect 41328 100 41384 400
rect 44016 100 44072 400
rect 46704 100 46760 400
rect 49056 100 49112 400
rect 51744 100 51800 400
rect 54432 100 54488 400
rect 57120 100 57176 400
rect 59472 100 59528 400
rect 62160 100 62216 400
rect 64848 100 64904 400
rect 67200 100 67256 400
rect 69888 100 69944 400
rect 72576 100 72632 400
rect 75264 100 75320 400
rect 77616 100 77672 400
rect 80304 100 80360 400
rect 82992 100 83048 400
rect 85680 100 85736 400
rect 88032 100 88088 400
rect 90720 100 90776 400
rect 93408 100 93464 400
rect 96096 100 96152 400
rect 98448 100 98504 400
rect 101136 100 101192 400
rect 103824 100 103880 400
rect 106176 100 106232 400
rect 108864 100 108920 400
rect 111552 100 111608 400
rect 114240 100 114296 400
rect 116592 100 116648 400
rect 119280 100 119336 400
rect 121968 100 122024 400
rect 124656 100 124712 400
rect 127008 100 127064 400
rect 129696 100 129752 400
rect 132384 100 132440 400
rect 134736 100 134792 400
rect 137424 100 137480 400
rect 140112 100 140168 400
rect 142800 100 142856 400
rect 145152 100 145208 400
rect 147840 100 147896 400
rect 150528 100 150584 400
rect 153216 100 153272 400
rect 155568 100 155624 400
rect 158256 100 158312 400
rect 160944 100 161000 400
rect 163296 100 163352 400
rect 165984 100 166040 400
rect 168672 100 168728 400
rect 171360 100 171416 400
rect 173712 100 173768 400
rect 176400 100 176456 400
rect 179088 100 179144 400
rect 181776 100 181832 400
rect 184128 100 184184 400
rect 186816 100 186872 400
rect 189504 100 189560 400
rect 192192 100 192248 400
rect 194544 100 194600 400
rect 197232 100 197288 400
rect 199920 100 199976 400
rect 202272 100 202328 400
rect 204960 100 205016 400
rect 207648 100 207704 400
rect 210336 100 210392 400
rect 212688 100 212744 400
rect 215376 100 215432 400
rect 218064 100 218120 400
rect 220752 100 220808 400
rect 223104 100 223160 400
rect 225792 100 225848 400
rect 228480 100 228536 400
rect 230832 100 230888 400
rect 233520 100 233576 400
rect 236208 100 236264 400
rect 238896 100 238952 400
rect 241248 100 241304 400
rect 243936 100 243992 400
rect 246624 100 246680 400
rect 249312 100 249368 400
<< obsm2 >>
rect 14 249930 249354 249970
rect 14 249570 1650 249930
rect 1766 249570 4338 249930
rect 4454 249570 7026 249930
rect 7142 249570 9378 249930
rect 9494 249570 12066 249930
rect 12182 249570 14754 249930
rect 14870 249570 17442 249930
rect 17558 249570 19794 249930
rect 19910 249570 22482 249930
rect 22598 249570 25170 249930
rect 25286 249570 27858 249930
rect 27974 249570 30210 249930
rect 30326 249570 32898 249930
rect 33014 249570 35586 249930
rect 35702 249570 38274 249930
rect 38390 249570 40626 249930
rect 40742 249570 43314 249930
rect 43430 249570 46002 249930
rect 46118 249570 48354 249930
rect 48470 249570 51042 249930
rect 51158 249570 53730 249930
rect 53846 249570 56418 249930
rect 56534 249570 58770 249930
rect 58886 249570 61458 249930
rect 61574 249570 64146 249930
rect 64262 249570 66834 249930
rect 66950 249570 69186 249930
rect 69302 249570 71874 249930
rect 71990 249570 74562 249930
rect 74678 249570 76914 249930
rect 77030 249570 79602 249930
rect 79718 249570 82290 249930
rect 82406 249570 84978 249930
rect 85094 249570 87330 249930
rect 87446 249570 90018 249930
rect 90134 249570 92706 249930
rect 92822 249570 95394 249930
rect 95510 249570 97746 249930
rect 97862 249570 100434 249930
rect 100550 249570 103122 249930
rect 103238 249570 105474 249930
rect 105590 249570 108162 249930
rect 108278 249570 110850 249930
rect 110966 249570 113538 249930
rect 113654 249570 115890 249930
rect 116006 249570 118578 249930
rect 118694 249570 121266 249930
rect 121382 249570 123954 249930
rect 124070 249570 126306 249930
rect 126422 249570 128994 249930
rect 129110 249570 131682 249930
rect 131798 249570 134370 249930
rect 134486 249570 136722 249930
rect 136838 249570 139410 249930
rect 139526 249570 142098 249930
rect 142214 249570 144450 249930
rect 144566 249570 147138 249930
rect 147254 249570 149826 249930
rect 149942 249570 152514 249930
rect 152630 249570 154866 249930
rect 154982 249570 157554 249930
rect 157670 249570 160242 249930
rect 160358 249570 162930 249930
rect 163046 249570 165282 249930
rect 165398 249570 167970 249930
rect 168086 249570 170658 249930
rect 170774 249570 173010 249930
rect 173126 249570 175698 249930
rect 175814 249570 178386 249930
rect 178502 249570 181074 249930
rect 181190 249570 183426 249930
rect 183542 249570 186114 249930
rect 186230 249570 188802 249930
rect 188918 249570 191490 249930
rect 191606 249570 193842 249930
rect 193958 249570 196530 249930
rect 196646 249570 199218 249930
rect 199334 249570 201570 249930
rect 201686 249570 204258 249930
rect 204374 249570 206946 249930
rect 207062 249570 209634 249930
rect 209750 249570 211986 249930
rect 212102 249570 214674 249930
rect 214790 249570 217362 249930
rect 217478 249570 220050 249930
rect 220166 249570 222402 249930
rect 222518 249570 225090 249930
rect 225206 249570 227778 249930
rect 227894 249570 230466 249930
rect 230582 249570 232818 249930
rect 232934 249570 235506 249930
rect 235622 249570 238194 249930
rect 238310 249570 240546 249930
rect 240662 249570 243234 249930
rect 243350 249570 245922 249930
rect 246038 249570 248610 249930
rect 248726 249570 249354 249930
rect 14 430 249354 249570
rect 86 350 2322 430
rect 2438 350 5010 430
rect 5126 350 7698 430
rect 7814 350 10050 430
rect 10166 350 12738 430
rect 12854 350 15426 430
rect 15542 350 18114 430
rect 18230 350 20466 430
rect 20582 350 23154 430
rect 23270 350 25842 430
rect 25958 350 28530 430
rect 28646 350 30882 430
rect 30998 350 33570 430
rect 33686 350 36258 430
rect 36374 350 38610 430
rect 38726 350 41298 430
rect 41414 350 43986 430
rect 44102 350 46674 430
rect 46790 350 49026 430
rect 49142 350 51714 430
rect 51830 350 54402 430
rect 54518 350 57090 430
rect 57206 350 59442 430
rect 59558 350 62130 430
rect 62246 350 64818 430
rect 64934 350 67170 430
rect 67286 350 69858 430
rect 69974 350 72546 430
rect 72662 350 75234 430
rect 75350 350 77586 430
rect 77702 350 80274 430
rect 80390 350 82962 430
rect 83078 350 85650 430
rect 85766 350 88002 430
rect 88118 350 90690 430
rect 90806 350 93378 430
rect 93494 350 96066 430
rect 96182 350 98418 430
rect 98534 350 101106 430
rect 101222 350 103794 430
rect 103910 350 106146 430
rect 106262 350 108834 430
rect 108950 350 111522 430
rect 111638 350 114210 430
rect 114326 350 116562 430
rect 116678 350 119250 430
rect 119366 350 121938 430
rect 122054 350 124626 430
rect 124742 350 126978 430
rect 127094 350 129666 430
rect 129782 350 132354 430
rect 132470 350 134706 430
rect 134822 350 137394 430
rect 137510 350 140082 430
rect 140198 350 142770 430
rect 142886 350 145122 430
rect 145238 350 147810 430
rect 147926 350 150498 430
rect 150614 350 153186 430
rect 153302 350 155538 430
rect 155654 350 158226 430
rect 158342 350 160914 430
rect 161030 350 163266 430
rect 163382 350 165954 430
rect 166070 350 168642 430
rect 168758 350 171330 430
rect 171446 350 173682 430
rect 173798 350 176370 430
rect 176486 350 179058 430
rect 179174 350 181746 430
rect 181862 350 184098 430
rect 184214 350 186786 430
rect 186902 350 189474 430
rect 189590 350 192162 430
rect 192278 350 194514 430
rect 194630 350 197202 430
rect 197318 350 199890 430
rect 200006 350 202242 430
rect 202358 350 204930 430
rect 205046 350 207618 430
rect 207734 350 210306 430
rect 210422 350 212658 430
rect 212774 350 215346 430
rect 215462 350 218034 430
rect 218150 350 220722 430
rect 220838 350 223074 430
rect 223190 350 225762 430
rect 225878 350 228450 430
rect 228566 350 230802 430
rect 230918 350 233490 430
rect 233606 350 236178 430
rect 236294 350 238866 430
rect 238982 350 241218 430
rect 241334 350 243906 430
rect 244022 350 246594 430
rect 246710 350 249282 430
<< metal3 >>
rect 100 249312 400 249368
rect 249600 248640 249900 248696
rect 100 246624 400 246680
rect 249600 245952 249900 246008
rect 100 243936 400 243992
rect 249600 243264 249900 243320
rect 100 241248 400 241304
rect 249600 240576 249900 240632
rect 100 238896 400 238952
rect 249600 238224 249900 238280
rect 100 236208 400 236264
rect 249600 235536 249900 235592
rect 100 233520 400 233576
rect 249600 232848 249900 232904
rect 100 230832 400 230888
rect 249600 230496 249900 230552
rect 100 228480 400 228536
rect 249600 227808 249900 227864
rect 100 225792 400 225848
rect 249600 225120 249900 225176
rect 100 223104 400 223160
rect 249600 222432 249900 222488
rect 100 220752 400 220808
rect 249600 220080 249900 220136
rect 100 218064 400 218120
rect 249600 217392 249900 217448
rect 100 215376 400 215432
rect 249600 214704 249900 214760
rect 100 212688 400 212744
rect 249600 212016 249900 212072
rect 100 210336 400 210392
rect 249600 209664 249900 209720
rect 100 207648 400 207704
rect 249600 206976 249900 207032
rect 100 204960 400 205016
rect 249600 204288 249900 204344
rect 100 202272 400 202328
rect 249600 201600 249900 201656
rect 100 199920 400 199976
rect 249600 199248 249900 199304
rect 100 197232 400 197288
rect 249600 196560 249900 196616
rect 100 194544 400 194600
rect 249600 193872 249900 193928
rect 100 192192 400 192248
rect 249600 191520 249900 191576
rect 100 189504 400 189560
rect 249600 188832 249900 188888
rect 100 186816 400 186872
rect 249600 186144 249900 186200
rect 100 184128 400 184184
rect 249600 183456 249900 183512
rect 100 181776 400 181832
rect 249600 181104 249900 181160
rect 100 179088 400 179144
rect 249600 178416 249900 178472
rect 100 176400 400 176456
rect 249600 175728 249900 175784
rect 100 173712 400 173768
rect 249600 173040 249900 173096
rect 100 171360 400 171416
rect 249600 170688 249900 170744
rect 100 168672 400 168728
rect 249600 168000 249900 168056
rect 100 165984 400 166040
rect 249600 165312 249900 165368
rect 100 163296 400 163352
rect 249600 162960 249900 163016
rect 100 160944 400 161000
rect 249600 160272 249900 160328
rect 100 158256 400 158312
rect 249600 157584 249900 157640
rect 100 155568 400 155624
rect 249600 154896 249900 154952
rect 100 153216 400 153272
rect 249600 152544 249900 152600
rect 100 150528 400 150584
rect 249600 149856 249900 149912
rect 100 147840 400 147896
rect 249600 147168 249900 147224
rect 100 145152 400 145208
rect 249600 144480 249900 144536
rect 100 142800 400 142856
rect 249600 142128 249900 142184
rect 100 140112 400 140168
rect 249600 139440 249900 139496
rect 100 137424 400 137480
rect 249600 136752 249900 136808
rect 100 134736 400 134792
rect 249600 134400 249900 134456
rect 100 132384 400 132440
rect 249600 131712 249900 131768
rect 100 129696 400 129752
rect 249600 129024 249900 129080
rect 100 127008 400 127064
rect 249600 126336 249900 126392
rect 100 124656 400 124712
rect 249600 123984 249900 124040
rect 100 121968 400 122024
rect 249600 121296 249900 121352
rect 100 119280 400 119336
rect 249600 118608 249900 118664
rect 100 116592 400 116648
rect 249600 115920 249900 115976
rect 100 114240 400 114296
rect 249600 113568 249900 113624
rect 100 111552 400 111608
rect 249600 110880 249900 110936
rect 100 108864 400 108920
rect 249600 108192 249900 108248
rect 100 106176 400 106232
rect 249600 105504 249900 105560
rect 100 103824 400 103880
rect 249600 103152 249900 103208
rect 100 101136 400 101192
rect 249600 100464 249900 100520
rect 100 98448 400 98504
rect 249600 97776 249900 97832
rect 100 96096 400 96152
rect 249600 95424 249900 95480
rect 100 93408 400 93464
rect 249600 92736 249900 92792
rect 100 90720 400 90776
rect 249600 90048 249900 90104
rect 100 88032 400 88088
rect 249600 87360 249900 87416
rect 100 85680 400 85736
rect 249600 85008 249900 85064
rect 100 82992 400 83048
rect 249600 82320 249900 82376
rect 100 80304 400 80360
rect 249600 79632 249900 79688
rect 100 77616 400 77672
rect 249600 76944 249900 77000
rect 100 75264 400 75320
rect 249600 74592 249900 74648
rect 100 72576 400 72632
rect 249600 71904 249900 71960
rect 100 69888 400 69944
rect 249600 69216 249900 69272
rect 100 67200 400 67256
rect 249600 66864 249900 66920
rect 100 64848 400 64904
rect 249600 64176 249900 64232
rect 100 62160 400 62216
rect 249600 61488 249900 61544
rect 100 59472 400 59528
rect 249600 58800 249900 58856
rect 100 57120 400 57176
rect 249600 56448 249900 56504
rect 100 54432 400 54488
rect 249600 53760 249900 53816
rect 100 51744 400 51800
rect 249600 51072 249900 51128
rect 100 49056 400 49112
rect 249600 48384 249900 48440
rect 100 46704 400 46760
rect 249600 46032 249900 46088
rect 100 44016 400 44072
rect 249600 43344 249900 43400
rect 100 41328 400 41384
rect 249600 40656 249900 40712
rect 100 38640 400 38696
rect 249600 38304 249900 38360
rect 100 36288 400 36344
rect 249600 35616 249900 35672
rect 100 33600 400 33656
rect 249600 32928 249900 32984
rect 100 30912 400 30968
rect 249600 30240 249900 30296
rect 100 28560 400 28616
rect 249600 27888 249900 27944
rect 100 25872 400 25928
rect 249600 25200 249900 25256
rect 100 23184 400 23240
rect 249600 22512 249900 22568
rect 100 20496 400 20552
rect 249600 19824 249900 19880
rect 100 18144 400 18200
rect 249600 17472 249900 17528
rect 100 15456 400 15512
rect 249600 14784 249900 14840
rect 100 12768 400 12824
rect 249600 12096 249900 12152
rect 100 10080 400 10136
rect 249600 9408 249900 9464
rect 100 7728 400 7784
rect 249600 7056 249900 7112
rect 100 5040 400 5096
rect 249600 4368 249900 4424
rect 100 2352 400 2408
rect 249600 1680 249900 1736
<< obsm3 >>
rect 9 249282 70 249354
rect 430 249282 249970 249354
rect 9 248726 249970 249282
rect 9 248610 249570 248726
rect 249930 248610 249970 248726
rect 9 246710 249970 248610
rect 9 246594 70 246710
rect 430 246594 249970 246710
rect 9 246038 249970 246594
rect 9 245922 249570 246038
rect 249930 245922 249970 246038
rect 9 244022 249970 245922
rect 9 243906 70 244022
rect 430 243906 249970 244022
rect 9 243350 249970 243906
rect 9 243234 249570 243350
rect 249930 243234 249970 243350
rect 9 241334 249970 243234
rect 9 241218 70 241334
rect 430 241218 249970 241334
rect 9 240662 249970 241218
rect 9 240546 249570 240662
rect 249930 240546 249970 240662
rect 9 238982 249970 240546
rect 9 238866 70 238982
rect 430 238866 249970 238982
rect 9 238310 249970 238866
rect 9 238194 249570 238310
rect 249930 238194 249970 238310
rect 9 236294 249970 238194
rect 9 236178 70 236294
rect 430 236178 249970 236294
rect 9 235622 249970 236178
rect 9 235506 249570 235622
rect 249930 235506 249970 235622
rect 9 233606 249970 235506
rect 9 233490 70 233606
rect 430 233490 249970 233606
rect 9 232934 249970 233490
rect 9 232818 249570 232934
rect 249930 232818 249970 232934
rect 9 230918 249970 232818
rect 9 230802 70 230918
rect 430 230802 249970 230918
rect 9 230582 249970 230802
rect 9 230466 249570 230582
rect 249930 230466 249970 230582
rect 9 228566 249970 230466
rect 9 228450 70 228566
rect 430 228450 249970 228566
rect 9 227894 249970 228450
rect 9 227778 249570 227894
rect 249930 227778 249970 227894
rect 9 225878 249970 227778
rect 9 225762 70 225878
rect 430 225762 249970 225878
rect 9 225206 249970 225762
rect 9 225090 249570 225206
rect 249930 225090 249970 225206
rect 9 223190 249970 225090
rect 9 223074 70 223190
rect 430 223074 249970 223190
rect 9 222518 249970 223074
rect 9 222402 249570 222518
rect 249930 222402 249970 222518
rect 9 220838 249970 222402
rect 9 220722 70 220838
rect 430 220722 249970 220838
rect 9 220166 249970 220722
rect 9 220050 249570 220166
rect 249930 220050 249970 220166
rect 9 218150 249970 220050
rect 9 218034 70 218150
rect 430 218034 249970 218150
rect 9 217478 249970 218034
rect 9 217362 249570 217478
rect 249930 217362 249970 217478
rect 9 215462 249970 217362
rect 9 215346 70 215462
rect 430 215346 249970 215462
rect 9 214790 249970 215346
rect 9 214674 249570 214790
rect 249930 214674 249970 214790
rect 9 212774 249970 214674
rect 9 212658 70 212774
rect 430 212658 249970 212774
rect 9 212102 249970 212658
rect 9 211986 249570 212102
rect 249930 211986 249970 212102
rect 9 210422 249970 211986
rect 9 210306 70 210422
rect 430 210306 249970 210422
rect 9 209750 249970 210306
rect 9 209634 249570 209750
rect 249930 209634 249970 209750
rect 9 207734 249970 209634
rect 9 207618 70 207734
rect 430 207618 249970 207734
rect 9 207062 249970 207618
rect 9 206946 249570 207062
rect 249930 206946 249970 207062
rect 9 205046 249970 206946
rect 9 204930 70 205046
rect 430 204930 249970 205046
rect 9 204374 249970 204930
rect 9 204258 249570 204374
rect 249930 204258 249970 204374
rect 9 202358 249970 204258
rect 9 202242 70 202358
rect 430 202242 249970 202358
rect 9 201686 249970 202242
rect 9 201570 249570 201686
rect 249930 201570 249970 201686
rect 9 200006 249970 201570
rect 9 199890 70 200006
rect 430 199890 249970 200006
rect 9 199334 249970 199890
rect 9 199218 249570 199334
rect 249930 199218 249970 199334
rect 9 197318 249970 199218
rect 9 197202 70 197318
rect 430 197202 249970 197318
rect 9 196646 249970 197202
rect 9 196530 249570 196646
rect 249930 196530 249970 196646
rect 9 194630 249970 196530
rect 9 194514 70 194630
rect 430 194514 249970 194630
rect 9 193958 249970 194514
rect 9 193842 249570 193958
rect 249930 193842 249970 193958
rect 9 192278 249970 193842
rect 9 192162 70 192278
rect 430 192162 249970 192278
rect 9 191606 249970 192162
rect 9 191490 249570 191606
rect 249930 191490 249970 191606
rect 9 189590 249970 191490
rect 9 189474 70 189590
rect 430 189474 249970 189590
rect 9 188918 249970 189474
rect 9 188802 249570 188918
rect 249930 188802 249970 188918
rect 9 186902 249970 188802
rect 9 186786 70 186902
rect 430 186786 249970 186902
rect 9 186230 249970 186786
rect 9 186114 249570 186230
rect 249930 186114 249970 186230
rect 9 184214 249970 186114
rect 9 184098 70 184214
rect 430 184098 249970 184214
rect 9 183542 249970 184098
rect 9 183426 249570 183542
rect 249930 183426 249970 183542
rect 9 181862 249970 183426
rect 9 181746 70 181862
rect 430 181746 249970 181862
rect 9 181190 249970 181746
rect 9 181074 249570 181190
rect 249930 181074 249970 181190
rect 9 179174 249970 181074
rect 9 179058 70 179174
rect 430 179058 249970 179174
rect 9 178502 249970 179058
rect 9 178386 249570 178502
rect 249930 178386 249970 178502
rect 9 176486 249970 178386
rect 9 176370 70 176486
rect 430 176370 249970 176486
rect 9 175814 249970 176370
rect 9 175698 249570 175814
rect 249930 175698 249970 175814
rect 9 173798 249970 175698
rect 9 173682 70 173798
rect 430 173682 249970 173798
rect 9 173126 249970 173682
rect 9 173010 249570 173126
rect 249930 173010 249970 173126
rect 9 171446 249970 173010
rect 9 171330 70 171446
rect 430 171330 249970 171446
rect 9 170774 249970 171330
rect 9 170658 249570 170774
rect 249930 170658 249970 170774
rect 9 168758 249970 170658
rect 9 168642 70 168758
rect 430 168642 249970 168758
rect 9 168086 249970 168642
rect 9 167970 249570 168086
rect 249930 167970 249970 168086
rect 9 166070 249970 167970
rect 9 165954 70 166070
rect 430 165954 249970 166070
rect 9 165398 249970 165954
rect 9 165282 249570 165398
rect 249930 165282 249970 165398
rect 9 163382 249970 165282
rect 9 163266 70 163382
rect 430 163266 249970 163382
rect 9 163046 249970 163266
rect 9 162930 249570 163046
rect 249930 162930 249970 163046
rect 9 161030 249970 162930
rect 9 160914 70 161030
rect 430 160914 249970 161030
rect 9 160358 249970 160914
rect 9 160242 249570 160358
rect 249930 160242 249970 160358
rect 9 158342 249970 160242
rect 9 158226 70 158342
rect 430 158226 249970 158342
rect 9 157670 249970 158226
rect 9 157554 249570 157670
rect 249930 157554 249970 157670
rect 9 155654 249970 157554
rect 9 155538 70 155654
rect 430 155538 249970 155654
rect 9 154982 249970 155538
rect 9 154866 249570 154982
rect 249930 154866 249970 154982
rect 9 153302 249970 154866
rect 9 153186 70 153302
rect 430 153186 249970 153302
rect 9 152630 249970 153186
rect 9 152514 249570 152630
rect 249930 152514 249970 152630
rect 9 150614 249970 152514
rect 9 150498 70 150614
rect 430 150498 249970 150614
rect 9 149942 249970 150498
rect 9 149826 249570 149942
rect 249930 149826 249970 149942
rect 9 147926 249970 149826
rect 9 147810 70 147926
rect 430 147810 249970 147926
rect 9 147254 249970 147810
rect 9 147138 249570 147254
rect 249930 147138 249970 147254
rect 9 145238 249970 147138
rect 9 145122 70 145238
rect 430 145122 249970 145238
rect 9 144566 249970 145122
rect 9 144450 249570 144566
rect 249930 144450 249970 144566
rect 9 142886 249970 144450
rect 9 142770 70 142886
rect 430 142770 249970 142886
rect 9 142214 249970 142770
rect 9 142098 249570 142214
rect 249930 142098 249970 142214
rect 9 140198 249970 142098
rect 9 140082 70 140198
rect 430 140082 249970 140198
rect 9 139526 249970 140082
rect 9 139410 249570 139526
rect 249930 139410 249970 139526
rect 9 137510 249970 139410
rect 9 137394 70 137510
rect 430 137394 249970 137510
rect 9 136838 249970 137394
rect 9 136722 249570 136838
rect 249930 136722 249970 136838
rect 9 134822 249970 136722
rect 9 134706 70 134822
rect 430 134706 249970 134822
rect 9 134486 249970 134706
rect 9 134370 249570 134486
rect 249930 134370 249970 134486
rect 9 132470 249970 134370
rect 9 132354 70 132470
rect 430 132354 249970 132470
rect 9 131798 249970 132354
rect 9 131682 249570 131798
rect 249930 131682 249970 131798
rect 9 129782 249970 131682
rect 9 129666 70 129782
rect 430 129666 249970 129782
rect 9 129110 249970 129666
rect 9 128994 249570 129110
rect 249930 128994 249970 129110
rect 9 127094 249970 128994
rect 9 126978 70 127094
rect 430 126978 249970 127094
rect 9 126422 249970 126978
rect 9 126306 249570 126422
rect 249930 126306 249970 126422
rect 9 124742 249970 126306
rect 9 124626 70 124742
rect 430 124626 249970 124742
rect 9 124070 249970 124626
rect 9 123954 249570 124070
rect 249930 123954 249970 124070
rect 9 122054 249970 123954
rect 9 121938 70 122054
rect 430 121938 249970 122054
rect 9 121382 249970 121938
rect 9 121266 249570 121382
rect 249930 121266 249970 121382
rect 9 119366 249970 121266
rect 9 119250 70 119366
rect 430 119250 249970 119366
rect 9 118694 249970 119250
rect 9 118578 249570 118694
rect 249930 118578 249970 118694
rect 9 116678 249970 118578
rect 9 116562 70 116678
rect 430 116562 249970 116678
rect 9 116006 249970 116562
rect 9 115890 249570 116006
rect 249930 115890 249970 116006
rect 9 114326 249970 115890
rect 9 114210 70 114326
rect 430 114210 249970 114326
rect 9 113654 249970 114210
rect 9 113538 249570 113654
rect 249930 113538 249970 113654
rect 9 111638 249970 113538
rect 9 111522 70 111638
rect 430 111522 249970 111638
rect 9 110966 249970 111522
rect 9 110850 249570 110966
rect 249930 110850 249970 110966
rect 9 108950 249970 110850
rect 9 108834 70 108950
rect 430 108834 249970 108950
rect 9 108278 249970 108834
rect 9 108162 249570 108278
rect 249930 108162 249970 108278
rect 9 106262 249970 108162
rect 9 106146 70 106262
rect 430 106146 249970 106262
rect 9 105590 249970 106146
rect 9 105474 249570 105590
rect 249930 105474 249970 105590
rect 9 103910 249970 105474
rect 9 103794 70 103910
rect 430 103794 249970 103910
rect 9 103238 249970 103794
rect 9 103122 249570 103238
rect 249930 103122 249970 103238
rect 9 101222 249970 103122
rect 9 101106 70 101222
rect 430 101106 249970 101222
rect 9 100550 249970 101106
rect 9 100434 249570 100550
rect 249930 100434 249970 100550
rect 9 98534 249970 100434
rect 9 98418 70 98534
rect 430 98418 249970 98534
rect 9 97862 249970 98418
rect 9 97746 249570 97862
rect 249930 97746 249970 97862
rect 9 96182 249970 97746
rect 9 96066 70 96182
rect 430 96066 249970 96182
rect 9 95510 249970 96066
rect 9 95394 249570 95510
rect 249930 95394 249970 95510
rect 9 93494 249970 95394
rect 9 93378 70 93494
rect 430 93378 249970 93494
rect 9 92822 249970 93378
rect 9 92706 249570 92822
rect 249930 92706 249970 92822
rect 9 90806 249970 92706
rect 9 90690 70 90806
rect 430 90690 249970 90806
rect 9 90134 249970 90690
rect 9 90018 249570 90134
rect 249930 90018 249970 90134
rect 9 88118 249970 90018
rect 9 88002 70 88118
rect 430 88002 249970 88118
rect 9 87446 249970 88002
rect 9 87330 249570 87446
rect 249930 87330 249970 87446
rect 9 85766 249970 87330
rect 9 85650 70 85766
rect 430 85650 249970 85766
rect 9 85094 249970 85650
rect 9 84978 249570 85094
rect 249930 84978 249970 85094
rect 9 83078 249970 84978
rect 9 82962 70 83078
rect 430 82962 249970 83078
rect 9 82406 249970 82962
rect 9 82290 249570 82406
rect 249930 82290 249970 82406
rect 9 80390 249970 82290
rect 9 80274 70 80390
rect 430 80274 249970 80390
rect 9 79718 249970 80274
rect 9 79602 249570 79718
rect 249930 79602 249970 79718
rect 9 77702 249970 79602
rect 9 77586 70 77702
rect 430 77586 249970 77702
rect 9 77030 249970 77586
rect 9 76914 249570 77030
rect 249930 76914 249970 77030
rect 9 75350 249970 76914
rect 9 75234 70 75350
rect 430 75234 249970 75350
rect 9 74678 249970 75234
rect 9 74562 249570 74678
rect 249930 74562 249970 74678
rect 9 72662 249970 74562
rect 9 72546 70 72662
rect 430 72546 249970 72662
rect 9 71990 249970 72546
rect 9 71874 249570 71990
rect 249930 71874 249970 71990
rect 9 69974 249970 71874
rect 9 69858 70 69974
rect 430 69858 249970 69974
rect 9 69302 249970 69858
rect 9 69186 249570 69302
rect 249930 69186 249970 69302
rect 9 67286 249970 69186
rect 9 67170 70 67286
rect 430 67170 249970 67286
rect 9 66950 249970 67170
rect 9 66834 249570 66950
rect 249930 66834 249970 66950
rect 9 64934 249970 66834
rect 9 64818 70 64934
rect 430 64818 249970 64934
rect 9 64262 249970 64818
rect 9 64146 249570 64262
rect 249930 64146 249970 64262
rect 9 62246 249970 64146
rect 9 62130 70 62246
rect 430 62130 249970 62246
rect 9 61574 249970 62130
rect 9 61458 249570 61574
rect 249930 61458 249970 61574
rect 9 59558 249970 61458
rect 9 59442 70 59558
rect 430 59442 249970 59558
rect 9 58886 249970 59442
rect 9 58770 249570 58886
rect 249930 58770 249970 58886
rect 9 57206 249970 58770
rect 9 57090 70 57206
rect 430 57090 249970 57206
rect 9 56534 249970 57090
rect 9 56418 249570 56534
rect 249930 56418 249970 56534
rect 9 54518 249970 56418
rect 9 54402 70 54518
rect 430 54402 249970 54518
rect 9 53846 249970 54402
rect 9 53730 249570 53846
rect 249930 53730 249970 53846
rect 9 51830 249970 53730
rect 9 51714 70 51830
rect 430 51714 249970 51830
rect 9 51158 249970 51714
rect 9 51042 249570 51158
rect 249930 51042 249970 51158
rect 9 49142 249970 51042
rect 9 49026 70 49142
rect 430 49026 249970 49142
rect 9 48470 249970 49026
rect 9 48354 249570 48470
rect 249930 48354 249970 48470
rect 9 46790 249970 48354
rect 9 46674 70 46790
rect 430 46674 249970 46790
rect 9 46118 249970 46674
rect 9 46002 249570 46118
rect 249930 46002 249970 46118
rect 9 44102 249970 46002
rect 9 43986 70 44102
rect 430 43986 249970 44102
rect 9 43430 249970 43986
rect 9 43314 249570 43430
rect 249930 43314 249970 43430
rect 9 41414 249970 43314
rect 9 41298 70 41414
rect 430 41298 249970 41414
rect 9 40742 249970 41298
rect 9 40626 249570 40742
rect 249930 40626 249970 40742
rect 9 38726 249970 40626
rect 9 38610 70 38726
rect 430 38610 249970 38726
rect 9 38390 249970 38610
rect 9 38274 249570 38390
rect 249930 38274 249970 38390
rect 9 36374 249970 38274
rect 9 36258 70 36374
rect 430 36258 249970 36374
rect 9 35702 249970 36258
rect 9 35586 249570 35702
rect 249930 35586 249970 35702
rect 9 33686 249970 35586
rect 9 33570 70 33686
rect 430 33570 249970 33686
rect 9 33014 249970 33570
rect 9 32898 249570 33014
rect 249930 32898 249970 33014
rect 9 30998 249970 32898
rect 9 30882 70 30998
rect 430 30882 249970 30998
rect 9 30326 249970 30882
rect 9 30210 249570 30326
rect 249930 30210 249970 30326
rect 9 28646 249970 30210
rect 9 28530 70 28646
rect 430 28530 249970 28646
rect 9 27974 249970 28530
rect 9 27858 249570 27974
rect 249930 27858 249970 27974
rect 9 25958 249970 27858
rect 9 25842 70 25958
rect 430 25842 249970 25958
rect 9 25286 249970 25842
rect 9 25170 249570 25286
rect 249930 25170 249970 25286
rect 9 23270 249970 25170
rect 9 23154 70 23270
rect 430 23154 249970 23270
rect 9 22598 249970 23154
rect 9 22482 249570 22598
rect 249930 22482 249970 22598
rect 9 20582 249970 22482
rect 9 20466 70 20582
rect 430 20466 249970 20582
rect 9 19910 249970 20466
rect 9 19794 249570 19910
rect 249930 19794 249970 19910
rect 9 18230 249970 19794
rect 9 18114 70 18230
rect 430 18114 249970 18230
rect 9 17558 249970 18114
rect 9 17442 249570 17558
rect 249930 17442 249970 17558
rect 9 15542 249970 17442
rect 9 15426 70 15542
rect 430 15426 249970 15542
rect 9 14870 249970 15426
rect 9 14754 249570 14870
rect 249930 14754 249970 14870
rect 9 12854 249970 14754
rect 9 12738 70 12854
rect 430 12738 249970 12854
rect 9 12182 249970 12738
rect 9 12066 249570 12182
rect 249930 12066 249970 12182
rect 9 10166 249970 12066
rect 9 10050 70 10166
rect 430 10050 249970 10166
rect 9 9494 249970 10050
rect 9 9378 249570 9494
rect 249930 9378 249970 9494
rect 9 7814 249970 9378
rect 9 7698 70 7814
rect 430 7698 249970 7814
rect 9 7142 249970 7698
rect 9 7026 249570 7142
rect 249930 7026 249970 7142
rect 9 5126 249970 7026
rect 9 5010 70 5126
rect 430 5010 249970 5126
rect 9 4454 249970 5010
rect 9 4338 249570 4454
rect 249930 4338 249970 4454
rect 9 2438 249970 4338
rect 9 2322 70 2438
rect 430 2322 249970 2438
rect 9 1766 249970 2322
rect 9 1650 249570 1766
rect 249930 1650 249970 1766
rect 9 574 249970 1650
<< metal4 >>
rect 2224 1538 2384 248166
rect 9904 1538 10064 248166
rect 17584 1538 17744 248166
rect 25264 1538 25424 248166
rect 32944 1538 33104 248166
rect 40624 1538 40784 248166
rect 48304 1538 48464 248166
rect 55984 1538 56144 248166
rect 63664 1538 63824 248166
rect 71344 1538 71504 248166
rect 79024 1538 79184 248166
rect 86704 1538 86864 248166
rect 94384 1538 94544 248166
rect 102064 1538 102224 248166
rect 109744 1538 109904 248166
rect 117424 1538 117584 248166
rect 125104 1538 125264 248166
rect 132784 1538 132944 248166
rect 140464 1538 140624 248166
rect 148144 1538 148304 248166
rect 155824 1538 155984 248166
rect 163504 1538 163664 248166
rect 171184 1538 171344 248166
rect 178864 1538 179024 248166
rect 186544 1538 186704 248166
rect 194224 1538 194384 248166
rect 201904 1538 202064 248166
rect 209584 1538 209744 248166
rect 217264 1538 217424 248166
rect 224944 1538 225104 248166
rect 232624 1538 232784 248166
rect 240304 1538 240464 248166
rect 247984 1538 248144 248166
<< obsm4 >>
rect 33502 2473 40594 247847
rect 40814 2473 48274 247847
rect 48494 2473 55954 247847
rect 56174 2473 63634 247847
rect 63854 2473 71314 247847
rect 71534 2473 78994 247847
rect 79214 2473 86674 247847
rect 86894 2473 94354 247847
rect 94574 2473 102034 247847
rect 102254 2473 109714 247847
rect 109934 2473 117394 247847
rect 117614 2473 125074 247847
rect 125294 2473 132754 247847
rect 132974 2473 140434 247847
rect 140654 2473 148114 247847
rect 148334 2473 155794 247847
rect 156014 2473 163474 247847
rect 163694 2473 171154 247847
rect 171374 2473 178834 247847
rect 179054 2473 186514 247847
rect 186734 2473 194194 247847
rect 194414 2473 201874 247847
rect 202094 2473 209554 247847
rect 209774 2473 217234 247847
rect 217454 2473 224914 247847
rect 225134 2473 232594 247847
rect 232814 2473 240274 247847
rect 240494 2473 247954 247847
rect 248174 2473 248850 247847
<< labels >>
rlabel metal3 s 100 103824 400 103880 6 clk
port 1 nsew signal input
rlabel metal2 s 232848 249600 232904 249900 6 key[0]
port 2 nsew signal input
rlabel metal3 s 100 59472 400 59528 6 key[100]
port 3 nsew signal input
rlabel metal2 s 204288 249600 204344 249900 6 key[101]
port 4 nsew signal input
rlabel metal3 s 100 15456 400 15512 6 key[102]
port 5 nsew signal input
rlabel metal3 s 100 150528 400 150584 6 key[103]
port 6 nsew signal input
rlabel metal3 s 100 137424 400 137480 6 key[104]
port 7 nsew signal input
rlabel metal3 s 249600 46032 249900 46088 6 key[105]
port 8 nsew signal input
rlabel metal3 s 100 218064 400 218120 6 key[106]
port 9 nsew signal input
rlabel metal2 s 100464 249600 100520 249900 6 key[107]
port 10 nsew signal input
rlabel metal2 s 85008 249600 85064 249900 6 key[108]
port 11 nsew signal input
rlabel metal2 s 170688 249600 170744 249900 6 key[109]
port 12 nsew signal input
rlabel metal3 s 249600 56448 249900 56504 6 key[10]
port 13 nsew signal input
rlabel metal2 s 222432 249600 222488 249900 6 key[110]
port 14 nsew signal input
rlabel metal3 s 100 160944 400 161000 6 key[111]
port 15 nsew signal input
rlabel metal2 s 132384 100 132440 400 6 key[112]
port 16 nsew signal input
rlabel metal3 s 249600 79632 249900 79688 6 key[113]
port 17 nsew signal input
rlabel metal2 s 240576 249600 240632 249900 6 key[114]
port 18 nsew signal input
rlabel metal3 s 100 199920 400 199976 6 key[115]
port 19 nsew signal input
rlabel metal3 s 100 64848 400 64904 6 key[116]
port 20 nsew signal input
rlabel metal3 s 249600 235536 249900 235592 6 key[117]
port 21 nsew signal input
rlabel metal3 s 249600 149856 249900 149912 6 key[118]
port 22 nsew signal input
rlabel metal2 s 225792 100 225848 400 6 key[119]
port 23 nsew signal input
rlabel metal2 s 193872 249600 193928 249900 6 key[11]
port 24 nsew signal input
rlabel metal2 s 158256 100 158312 400 6 key[120]
port 25 nsew signal input
rlabel metal3 s 100 243936 400 243992 6 key[121]
port 26 nsew signal input
rlabel metal2 s 95424 249600 95480 249900 6 key[122]
port 27 nsew signal input
rlabel metal3 s 249600 212016 249900 212072 6 key[123]
port 28 nsew signal input
rlabel metal3 s 249600 90048 249900 90104 6 key[124]
port 29 nsew signal input
rlabel metal3 s 100 238896 400 238952 6 key[125]
port 30 nsew signal input
rlabel metal2 s 186144 249600 186200 249900 6 key[126]
port 31 nsew signal input
rlabel metal3 s 249600 181104 249900 181160 6 key[127]
port 32 nsew signal input
rlabel metal2 s 57120 100 57176 400 6 key[12]
port 33 nsew signal input
rlabel metal3 s 249600 131712 249900 131768 6 key[13]
port 34 nsew signal input
rlabel metal2 s 15456 100 15512 400 6 key[14]
port 35 nsew signal input
rlabel metal2 s 243936 100 243992 400 6 key[15]
port 36 nsew signal input
rlabel metal2 s 153216 100 153272 400 6 key[16]
port 37 nsew signal input
rlabel metal3 s 100 77616 400 77672 6 key[17]
port 38 nsew signal input
rlabel metal3 s 100 80304 400 80360 6 key[18]
port 39 nsew signal input
rlabel metal3 s 249600 58800 249900 58856 6 key[19]
port 40 nsew signal input
rlabel metal3 s 249600 232848 249900 232904 6 key[1]
port 41 nsew signal input
rlabel metal2 s 220752 100 220808 400 6 key[20]
port 42 nsew signal input
rlabel metal3 s 249600 168000 249900 168056 6 key[21]
port 43 nsew signal input
rlabel metal3 s 249600 248640 249900 248696 6 key[22]
port 44 nsew signal input
rlabel metal2 s 163296 100 163352 400 6 key[23]
port 45 nsew signal input
rlabel metal3 s 100 20496 400 20552 6 key[24]
port 46 nsew signal input
rlabel metal2 s 61488 249600 61544 249900 6 key[25]
port 47 nsew signal input
rlabel metal2 s 56448 249600 56504 249900 6 key[26]
port 48 nsew signal input
rlabel metal2 s 126336 249600 126392 249900 6 key[27]
port 49 nsew signal input
rlabel metal3 s 100 186816 400 186872 6 key[28]
port 50 nsew signal input
rlabel metal2 s 23184 100 23240 400 6 key[29]
port 51 nsew signal input
rlabel metal3 s 249600 199248 249900 199304 6 key[2]
port 52 nsew signal input
rlabel metal3 s 249600 121296 249900 121352 6 key[30]
port 53 nsew signal input
rlabel metal2 s 9408 249600 9464 249900 6 key[31]
port 54 nsew signal input
rlabel metal2 s 233520 100 233576 400 6 key[32]
port 55 nsew signal input
rlabel metal3 s 249600 32928 249900 32984 6 key[33]
port 56 nsew signal input
rlabel metal3 s 249600 154896 249900 154952 6 key[34]
port 57 nsew signal input
rlabel metal3 s 100 38640 400 38696 6 key[35]
port 58 nsew signal input
rlabel metal3 s 249600 245952 249900 246008 6 key[36]
port 59 nsew signal input
rlabel metal3 s 249600 110880 249900 110936 6 key[37]
port 60 nsew signal input
rlabel metal3 s 249600 222432 249900 222488 6 key[38]
port 61 nsew signal input
rlabel metal3 s 100 181776 400 181832 6 key[39]
port 62 nsew signal input
rlabel metal2 s 160272 249600 160328 249900 6 key[3]
port 63 nsew signal input
rlabel metal3 s 100 194544 400 194600 6 key[40]
port 64 nsew signal input
rlabel metal2 s 59472 100 59528 400 6 key[41]
port 65 nsew signal input
rlabel metal2 s 215376 100 215432 400 6 key[42]
port 66 nsew signal input
rlabel metal2 s 121296 249600 121352 249900 6 key[43]
port 67 nsew signal input
rlabel metal2 s 176400 100 176456 400 6 key[44]
port 68 nsew signal input
rlabel metal2 s 199248 249600 199304 249900 6 key[45]
port 69 nsew signal input
rlabel metal2 s 241248 100 241304 400 6 key[46]
port 70 nsew signal input
rlabel metal2 s 140112 100 140168 400 6 key[47]
port 71 nsew signal input
rlabel metal2 s 144480 249600 144536 249900 6 key[48]
port 72 nsew signal input
rlabel metal2 s 127008 100 127064 400 6 key[49]
port 73 nsew signal input
rlabel metal3 s 249600 201600 249900 201656 6 key[4]
port 74 nsew signal input
rlabel metal2 s 105504 249600 105560 249900 6 key[50]
port 75 nsew signal input
rlabel metal3 s 249600 129024 249900 129080 6 key[51]
port 76 nsew signal input
rlabel metal2 s 194544 100 194600 400 6 key[52]
port 77 nsew signal input
rlabel metal3 s 249600 188832 249900 188888 6 key[53]
port 78 nsew signal input
rlabel metal3 s 249600 186144 249900 186200 6 key[54]
port 79 nsew signal input
rlabel metal2 s 108864 100 108920 400 6 key[55]
port 80 nsew signal input
rlabel metal2 s 28560 100 28616 400 6 key[56]
port 81 nsew signal input
rlabel metal3 s 100 163296 400 163352 6 key[57]
port 82 nsew signal input
rlabel metal3 s 249600 48384 249900 48440 6 key[58]
port 83 nsew signal input
rlabel metal2 s 48384 249600 48440 249900 6 key[59]
port 84 nsew signal input
rlabel metal2 s 199920 100 199976 400 6 key[5]
port 85 nsew signal input
rlabel metal3 s 249600 4368 249900 4424 6 key[60]
port 86 nsew signal input
rlabel metal2 s 4368 249600 4424 249900 6 key[61]
port 87 nsew signal input
rlabel metal3 s 100 93408 400 93464 6 key[62]
port 88 nsew signal input
rlabel metal3 s 249600 238224 249900 238280 6 key[63]
port 89 nsew signal input
rlabel metal2 s 93408 100 93464 400 6 key[64]
port 90 nsew signal input
rlabel metal2 s 116592 100 116648 400 6 key[65]
port 91 nsew signal input
rlabel metal2 s 40656 249600 40712 249900 6 key[66]
port 92 nsew signal input
rlabel metal3 s 249600 217392 249900 217448 6 key[67]
port 93 nsew signal input
rlabel metal2 s 64176 249600 64232 249900 6 key[68]
port 94 nsew signal input
rlabel metal2 s 14784 249600 14840 249900 6 key[69]
port 95 nsew signal input
rlabel metal3 s 100 189504 400 189560 6 key[6]
port 96 nsew signal input
rlabel metal2 s 35616 249600 35672 249900 6 key[70]
port 97 nsew signal input
rlabel metal3 s 249600 61488 249900 61544 6 key[71]
port 98 nsew signal input
rlabel metal2 s 75264 100 75320 400 6 key[72]
port 99 nsew signal input
rlabel metal2 s 113568 249600 113624 249900 6 key[73]
port 100 nsew signal input
rlabel metal3 s 100 62160 400 62216 6 key[74]
port 101 nsew signal input
rlabel metal2 s 123984 249600 124040 249900 6 key[75]
port 102 nsew signal input
rlabel metal3 s 249600 25200 249900 25256 6 key[76]
port 103 nsew signal input
rlabel metal2 s 64848 100 64904 400 6 key[77]
port 104 nsew signal input
rlabel metal2 s 147168 249600 147224 249900 6 key[78]
port 105 nsew signal input
rlabel metal3 s 249600 170688 249900 170744 6 key[79]
port 106 nsew signal input
rlabel metal3 s 249600 17472 249900 17528 6 key[7]
port 107 nsew signal input
rlabel metal2 s 248640 249600 248696 249900 6 key[80]
port 108 nsew signal input
rlabel metal3 s 100 142800 400 142856 6 key[81]
port 109 nsew signal input
rlabel metal2 s 149856 249600 149912 249900 6 key[82]
port 110 nsew signal input
rlabel metal2 s 217392 249600 217448 249900 6 key[83]
port 111 nsew signal input
rlabel metal3 s 249600 206976 249900 207032 6 key[84]
port 112 nsew signal input
rlabel metal3 s 100 28560 400 28616 6 key[85]
port 113 nsew signal input
rlabel metal3 s 249600 204288 249900 204344 6 key[86]
port 114 nsew signal input
rlabel metal3 s 100 108864 400 108920 6 key[87]
port 115 nsew signal input
rlabel metal2 s 49056 100 49112 400 6 key[88]
port 116 nsew signal input
rlabel metal2 s 25200 249600 25256 249900 6 key[89]
port 117 nsew signal input
rlabel metal3 s 100 173712 400 173768 6 key[8]
port 118 nsew signal input
rlabel metal2 s 103824 100 103880 400 6 key[90]
port 119 nsew signal input
rlabel metal2 s 82992 100 83048 400 6 key[91]
port 120 nsew signal input
rlabel metal2 s 36288 100 36344 400 6 key[92]
port 121 nsew signal input
rlabel metal2 s 218064 100 218120 400 6 key[93]
port 122 nsew signal input
rlabel metal2 s 69888 100 69944 400 6 key[94]
port 123 nsew signal input
rlabel metal3 s 100 249312 400 249368 6 key[95]
port 124 nsew signal input
rlabel metal3 s 100 176400 400 176456 6 key[96]
port 125 nsew signal input
rlabel metal2 s 74592 249600 74648 249900 6 key[97]
port 126 nsew signal input
rlabel metal3 s 100 75264 400 75320 6 key[98]
port 127 nsew signal input
rlabel metal2 s 115920 249600 115976 249900 6 key[99]
port 128 nsew signal input
rlabel metal3 s 249600 95424 249900 95480 6 key[9]
port 129 nsew signal input
rlabel metal2 s 101136 100 101192 400 6 out[0]
port 130 nsew signal output
rlabel metal3 s 249600 40656 249900 40712 6 out[100]
port 131 nsew signal output
rlabel metal2 s 1680 249600 1736 249900 6 out[101]
port 132 nsew signal output
rlabel metal3 s 249600 30240 249900 30296 6 out[102]
port 133 nsew signal output
rlabel metal3 s 100 72576 400 72632 6 out[103]
port 134 nsew signal output
rlabel metal3 s 100 5040 400 5096 6 out[104]
port 135 nsew signal output
rlabel metal2 s 228480 100 228536 400 6 out[105]
port 136 nsew signal output
rlabel metal2 s 80304 100 80360 400 6 out[106]
port 137 nsew signal output
rlabel metal2 s 209664 249600 209720 249900 6 out[107]
port 138 nsew signal output
rlabel metal3 s 100 153216 400 153272 6 out[108]
port 139 nsew signal output
rlabel metal2 s 19824 249600 19880 249900 6 out[109]
port 140 nsew signal output
rlabel metal2 s 114240 100 114296 400 6 out[10]
port 141 nsew signal output
rlabel metal3 s 100 236208 400 236264 6 out[110]
port 142 nsew signal output
rlabel metal2 s 139440 249600 139496 249900 6 out[111]
port 143 nsew signal output
rlabel metal2 s 152544 249600 152600 249900 6 out[112]
port 144 nsew signal output
rlabel metal3 s 249600 53760 249900 53816 6 out[113]
port 145 nsew signal output
rlabel metal3 s 249600 225120 249900 225176 6 out[114]
port 146 nsew signal output
rlabel metal2 s 204960 100 205016 400 6 out[115]
port 147 nsew signal output
rlabel metal3 s 249600 87360 249900 87416 6 out[116]
port 148 nsew signal output
rlabel metal3 s 249600 92736 249900 92792 6 out[117]
port 149 nsew signal output
rlabel metal2 s 160944 100 161000 400 6 out[118]
port 150 nsew signal output
rlabel metal2 s 72576 100 72632 400 6 out[119]
port 151 nsew signal output
rlabel metal2 s 85680 100 85736 400 6 out[11]
port 152 nsew signal output
rlabel metal3 s 249600 66864 249900 66920 6 out[120]
port 153 nsew signal output
rlabel metal3 s 249600 196560 249900 196616 6 out[121]
port 154 nsew signal output
rlabel metal3 s 100 179088 400 179144 6 out[122]
port 155 nsew signal output
rlabel metal2 s 41328 100 41384 400 6 out[123]
port 156 nsew signal output
rlabel metal3 s 249600 162960 249900 163016 6 out[124]
port 157 nsew signal output
rlabel metal3 s 100 155568 400 155624 6 out[125]
port 158 nsew signal output
rlabel metal3 s 249600 82320 249900 82376 6 out[126]
port 159 nsew signal output
rlabel metal2 s 12096 249600 12152 249900 6 out[127]
port 160 nsew signal output
rlabel metal3 s 249600 136752 249900 136808 6 out[12]
port 161 nsew signal output
rlabel metal2 s 154896 249600 154952 249900 6 out[13]
port 162 nsew signal output
rlabel metal3 s 100 18144 400 18200 6 out[14]
port 163 nsew signal output
rlabel metal3 s 249600 43344 249900 43400 6 out[15]
port 164 nsew signal output
rlabel metal2 s 134400 249600 134456 249900 6 out[16]
port 165 nsew signal output
rlabel metal3 s 100 44016 400 44072 6 out[17]
port 166 nsew signal output
rlabel metal2 s 53760 249600 53816 249900 6 out[18]
port 167 nsew signal output
rlabel metal3 s 249600 160272 249900 160328 6 out[19]
port 168 nsew signal output
rlabel metal2 s 98448 100 98504 400 6 out[1]
port 169 nsew signal output
rlabel metal2 s 88032 100 88088 400 6 out[20]
port 170 nsew signal output
rlabel metal3 s 249600 85008 249900 85064 6 out[21]
port 171 nsew signal output
rlabel metal2 s 79632 249600 79688 249900 6 out[22]
port 172 nsew signal output
rlabel metal2 s 38304 249600 38360 249900 6 out[23]
port 173 nsew signal output
rlabel metal3 s 249600 22512 249900 22568 6 out[24]
port 174 nsew signal output
rlabel metal2 s 111552 100 111608 400 6 out[25]
port 175 nsew signal output
rlabel metal2 s 220080 249600 220136 249900 6 out[26]
port 176 nsew signal output
rlabel metal3 s 249600 165312 249900 165368 6 out[27]
port 177 nsew signal output
rlabel metal3 s 100 41328 400 41384 6 out[28]
port 178 nsew signal output
rlabel metal3 s 100 241248 400 241304 6 out[29]
port 179 nsew signal output
rlabel metal3 s 100 101136 400 101192 6 out[2]
port 180 nsew signal output
rlabel metal2 s 145152 100 145208 400 6 out[30]
port 181 nsew signal output
rlabel metal2 s 58800 249600 58856 249900 6 out[31]
port 182 nsew signal output
rlabel metal2 s 212016 249600 212072 249900 6 out[32]
port 183 nsew signal output
rlabel metal3 s 249600 175728 249900 175784 6 out[33]
port 184 nsew signal output
rlabel metal2 s 12768 100 12824 400 6 out[34]
port 185 nsew signal output
rlabel metal3 s 100 210336 400 210392 6 out[35]
port 186 nsew signal output
rlabel metal2 s 17472 249600 17528 249900 6 out[36]
port 187 nsew signal output
rlabel metal2 s 157584 249600 157640 249900 6 out[37]
port 188 nsew signal output
rlabel metal3 s 100 192192 400 192248 6 out[38]
port 189 nsew signal output
rlabel metal3 s 100 33600 400 33656 6 out[39]
port 190 nsew signal output
rlabel metal2 s 210336 100 210392 400 6 out[3]
port 191 nsew signal output
rlabel metal3 s 249600 103152 249900 103208 6 out[40]
port 192 nsew signal output
rlabel metal3 s 249600 9408 249900 9464 6 out[41]
port 193 nsew signal output
rlabel metal3 s 100 7728 400 7784 6 out[42]
port 194 nsew signal output
rlabel metal2 s 110880 249600 110936 249900 6 out[43]
port 195 nsew signal output
rlabel metal2 s 129696 100 129752 400 6 out[44]
port 196 nsew signal output
rlabel metal3 s 100 246624 400 246680 6 out[45]
port 197 nsew signal output
rlabel metal2 s 119280 100 119336 400 6 out[46]
port 198 nsew signal output
rlabel metal3 s 249600 38304 249900 38360 6 out[47]
port 199 nsew signal output
rlabel metal2 s 225120 249600 225176 249900 6 out[48]
port 200 nsew signal output
rlabel metal3 s 100 49056 400 49112 6 out[49]
port 201 nsew signal output
rlabel metal2 s 142128 249600 142184 249900 6 out[4]
port 202 nsew signal output
rlabel metal3 s 100 88032 400 88088 6 out[50]
port 203 nsew signal output
rlabel metal2 s 235536 249600 235592 249900 6 out[51]
port 204 nsew signal output
rlabel metal2 s 43344 249600 43400 249900 6 out[52]
port 205 nsew signal output
rlabel metal3 s 100 67200 400 67256 6 out[53]
port 206 nsew signal output
rlabel metal3 s 249600 1680 249900 1736 6 out[54]
port 207 nsew signal output
rlabel metal3 s 100 228480 400 228536 6 out[55]
port 208 nsew signal output
rlabel metal3 s 100 212688 400 212744 6 out[56]
port 209 nsew signal output
rlabel metal2 s 147840 100 147896 400 6 out[57]
port 210 nsew signal output
rlabel metal3 s 249600 97776 249900 97832 6 out[58]
port 211 nsew signal output
rlabel metal3 s 249600 74592 249900 74648 6 out[59]
port 212 nsew signal output
rlabel metal2 s 87360 249600 87416 249900 6 out[5]
port 213 nsew signal output
rlabel metal3 s 249600 118608 249900 118664 6 out[60]
port 214 nsew signal output
rlabel metal2 s 179088 100 179144 400 6 out[61]
port 215 nsew signal output
rlabel metal3 s 100 2352 400 2408 6 out[62]
port 216 nsew signal output
rlabel metal2 s 173712 100 173768 400 6 out[63]
port 217 nsew signal output
rlabel metal2 s 207648 100 207704 400 6 out[64]
port 218 nsew signal output
rlabel metal2 s 33600 100 33656 400 6 out[65]
port 219 nsew signal output
rlabel metal3 s 100 168672 400 168728 6 out[66]
port 220 nsew signal output
rlabel metal2 s 189504 100 189560 400 6 out[67]
port 221 nsew signal output
rlabel metal3 s 100 116592 400 116648 6 out[68]
port 222 nsew signal output
rlabel metal3 s 100 184128 400 184184 6 out[69]
port 223 nsew signal output
rlabel metal3 s 249600 243264 249900 243320 6 out[6]
port 224 nsew signal output
rlabel metal3 s 100 51744 400 51800 6 out[70]
port 225 nsew signal output
rlabel metal3 s 100 134736 400 134792 6 out[71]
port 226 nsew signal output
rlabel metal2 s 67200 100 67256 400 6 out[72]
port 227 nsew signal output
rlabel metal3 s 249600 134400 249900 134456 6 out[73]
port 228 nsew signal output
rlabel metal2 s 212688 100 212744 400 6 out[74]
port 229 nsew signal output
rlabel metal2 s 196560 249600 196616 249900 6 out[75]
port 230 nsew signal output
rlabel metal2 s 44016 100 44072 400 6 out[76]
port 231 nsew signal output
rlabel metal2 s 51072 249600 51128 249900 6 out[77]
port 232 nsew signal output
rlabel metal3 s 249600 214704 249900 214760 6 out[78]
port 233 nsew signal output
rlabel metal3 s 100 90720 400 90776 6 out[79]
port 234 nsew signal output
rlabel metal3 s 249600 193872 249900 193928 6 out[7]
port 235 nsew signal output
rlabel metal2 s 136752 249600 136808 249900 6 out[80]
port 236 nsew signal output
rlabel metal3 s 100 25872 400 25928 6 out[81]
port 237 nsew signal output
rlabel metal3 s 100 111552 400 111608 6 out[82]
port 238 nsew signal output
rlabel metal3 s 100 147840 400 147896 6 out[83]
port 239 nsew signal output
rlabel metal2 s 108192 249600 108248 249900 6 out[84]
port 240 nsew signal output
rlabel metal2 s 2352 100 2408 400 6 out[85]
port 241 nsew signal output
rlabel metal2 s 69216 249600 69272 249900 6 out[86]
port 242 nsew signal output
rlabel metal2 s 124656 100 124712 400 6 out[87]
port 243 nsew signal output
rlabel metal2 s 249312 100 249368 400 6 out[88]
port 244 nsew signal output
rlabel metal3 s 249600 240576 249900 240632 6 out[89]
port 245 nsew signal output
rlabel metal3 s 249600 19824 249900 19880 6 out[8]
port 246 nsew signal output
rlabel metal2 s 118608 249600 118664 249900 6 out[90]
port 247 nsew signal output
rlabel metal2 s 7728 100 7784 400 6 out[91]
port 248 nsew signal output
rlabel metal2 s 46704 100 46760 400 6 out[92]
port 249 nsew signal output
rlabel metal2 s 106176 100 106232 400 6 out[93]
port 250 nsew signal output
rlabel metal2 s 227808 249600 227864 249900 6 out[94]
port 251 nsew signal output
rlabel metal3 s 100 202272 400 202328 6 out[95]
port 252 nsew signal output
rlabel metal2 s 90720 100 90776 400 6 out[96]
port 253 nsew signal output
rlabel metal3 s 100 10080 400 10136 6 out[97]
port 254 nsew signal output
rlabel metal3 s 249600 108192 249900 108248 6 out[98]
port 255 nsew signal output
rlabel metal3 s 100 225792 400 225848 6 out[99]
port 256 nsew signal output
rlabel metal2 s 186816 100 186872 400 6 out[9]
port 257 nsew signal output
rlabel metal3 s 100 12768 400 12824 6 state[0]
port 258 nsew signal input
rlabel metal2 s 238896 100 238952 400 6 state[100]
port 259 nsew signal input
rlabel metal3 s 249600 144480 249900 144536 6 state[101]
port 260 nsew signal input
rlabel metal2 s 188832 249600 188888 249900 6 state[102]
port 261 nsew signal input
rlabel metal3 s 249600 115920 249900 115976 6 state[103]
port 262 nsew signal input
rlabel metal3 s 100 197232 400 197288 6 state[104]
port 263 nsew signal input
rlabel metal3 s 100 145152 400 145208 6 state[105]
port 264 nsew signal input
rlabel metal3 s 249600 14784 249900 14840 6 state[106]
port 265 nsew signal input
rlabel metal2 s 168000 249600 168056 249900 6 state[107]
port 266 nsew signal input
rlabel metal2 s 223104 100 223160 400 6 state[108]
port 267 nsew signal input
rlabel metal2 s 30240 249600 30296 249900 6 state[109]
port 268 nsew signal input
rlabel metal2 s 30912 100 30968 400 6 state[10]
port 269 nsew signal input
rlabel metal3 s 249600 113568 249900 113624 6 state[110]
port 270 nsew signal input
rlabel metal2 s 7056 249600 7112 249900 6 state[111]
port 271 nsew signal input
rlabel metal3 s 249600 152544 249900 152600 6 state[112]
port 272 nsew signal input
rlabel metal2 s 62160 100 62216 400 6 state[113]
port 273 nsew signal input
rlabel metal2 s 230832 100 230888 400 6 state[114]
port 274 nsew signal input
rlabel metal2 s 92736 249600 92792 249900 6 state[115]
port 275 nsew signal input
rlabel metal2 s 230496 249600 230552 249900 6 state[116]
port 276 nsew signal input
rlabel metal3 s 249600 178416 249900 178472 6 state[117]
port 277 nsew signal input
rlabel metal2 s 82320 249600 82376 249900 6 state[118]
port 278 nsew signal input
rlabel metal2 s 103152 249600 103208 249900 6 state[119]
port 279 nsew signal input
rlabel metal3 s 249600 35616 249900 35672 6 state[11]
port 280 nsew signal input
rlabel metal3 s 100 132384 400 132440 6 state[120]
port 281 nsew signal input
rlabel metal3 s 100 119280 400 119336 6 state[121]
port 282 nsew signal input
rlabel metal2 s 181104 249600 181160 249900 6 state[122]
port 283 nsew signal input
rlabel metal2 s 129024 249600 129080 249900 6 state[123]
port 284 nsew signal input
rlabel metal2 s 32928 249600 32984 249900 6 state[124]
port 285 nsew signal input
rlabel metal3 s 100 98448 400 98504 6 state[125]
port 286 nsew signal input
rlabel metal3 s 100 233520 400 233576 6 state[126]
port 287 nsew signal input
rlabel metal3 s 249600 173040 249900 173096 6 state[127]
port 288 nsew signal input
rlabel metal3 s 249600 157584 249900 157640 6 state[12]
port 289 nsew signal input
rlabel metal2 s 155568 100 155624 400 6 state[13]
port 290 nsew signal input
rlabel metal3 s 249600 142128 249900 142184 6 state[14]
port 291 nsew signal input
rlabel metal3 s 100 121968 400 122024 6 state[15]
port 292 nsew signal input
rlabel metal2 s 236208 100 236264 400 6 state[16]
port 293 nsew signal input
rlabel metal2 s 173040 249600 173096 249900 6 state[17]
port 294 nsew signal input
rlabel metal2 s 243264 249600 243320 249900 6 state[18]
port 295 nsew signal input
rlabel metal2 s 137424 100 137480 400 6 state[19]
port 296 nsew signal input
rlabel metal3 s 100 69888 400 69944 6 state[1]
port 297 nsew signal input
rlabel metal3 s 249600 51072 249900 51128 6 state[20]
port 298 nsew signal input
rlabel metal2 s 46032 249600 46088 249900 6 state[21]
port 299 nsew signal input
rlabel metal3 s 100 46704 400 46760 6 state[22]
port 300 nsew signal input
rlabel metal2 s 25872 100 25928 400 6 state[23]
port 301 nsew signal input
rlabel metal2 s 97776 249600 97832 249900 6 state[24]
port 302 nsew signal input
rlabel metal3 s 100 96096 400 96152 6 state[25]
port 303 nsew signal input
rlabel metal3 s 249600 230496 249900 230552 6 state[26]
port 304 nsew signal input
rlabel metal3 s 100 30912 400 30968 6 state[27]
port 305 nsew signal input
rlabel metal2 s 206976 249600 207032 249900 6 state[28]
port 306 nsew signal input
rlabel metal3 s 249600 100464 249900 100520 6 state[29]
port 307 nsew signal input
rlabel metal2 s 192192 100 192248 400 6 state[2]
port 308 nsew signal input
rlabel metal3 s 100 106176 400 106232 6 state[30]
port 309 nsew signal input
rlabel metal2 s 184128 100 184184 400 6 state[31]
port 310 nsew signal input
rlabel metal3 s 100 129696 400 129752 6 state[32]
port 311 nsew signal input
rlabel metal3 s 100 171360 400 171416 6 state[33]
port 312 nsew signal input
rlabel metal2 s 246624 100 246680 400 6 state[34]
port 313 nsew signal input
rlabel metal3 s 249600 64176 249900 64232 6 state[35]
port 314 nsew signal input
rlabel metal2 s 90048 249600 90104 249900 6 state[36]
port 315 nsew signal input
rlabel metal3 s 249600 209664 249900 209720 6 state[37]
port 316 nsew signal input
rlabel metal3 s 100 204960 400 205016 6 state[38]
port 317 nsew signal input
rlabel metal3 s 100 223104 400 223160 6 state[39]
port 318 nsew signal input
rlabel metal3 s 100 215376 400 215432 6 state[3]
port 319 nsew signal input
rlabel metal2 s 10080 100 10136 400 6 state[40]
port 320 nsew signal input
rlabel metal3 s 100 57120 400 57176 6 state[41]
port 321 nsew signal input
rlabel metal3 s 249600 126336 249900 126392 6 state[42]
port 322 nsew signal input
rlabel metal2 s 142800 100 142856 400 6 state[43]
port 323 nsew signal input
rlabel metal2 s 178416 249600 178472 249900 6 state[44]
port 324 nsew signal input
rlabel metal2 s 238224 249600 238280 249900 6 state[45]
port 325 nsew signal input
rlabel metal2 s 22512 249600 22568 249900 6 state[46]
port 326 nsew signal input
rlabel metal3 s 100 114240 400 114296 6 state[47]
port 327 nsew signal input
rlabel metal3 s 100 127008 400 127064 6 state[48]
port 328 nsew signal input
rlabel metal2 s 245952 249600 246008 249900 6 state[49]
port 329 nsew signal input
rlabel metal3 s 100 158256 400 158312 6 state[4]
port 330 nsew signal input
rlabel metal3 s 100 36288 400 36344 6 state[50]
port 331 nsew signal input
rlabel metal3 s 249600 76944 249900 77000 6 state[51]
port 332 nsew signal input
rlabel metal2 s 171360 100 171416 400 6 state[52]
port 333 nsew signal input
rlabel metal2 s 214704 249600 214760 249900 6 state[53]
port 334 nsew signal input
rlabel metal2 s 66864 249600 66920 249900 6 state[54]
port 335 nsew signal input
rlabel metal2 s 77616 100 77672 400 6 state[55]
port 336 nsew signal input
rlabel metal3 s 249600 147168 249900 147224 6 state[56]
port 337 nsew signal input
rlabel metal2 s 202272 100 202328 400 6 state[57]
port 338 nsew signal input
rlabel metal3 s 249600 71904 249900 71960 6 state[58]
port 339 nsew signal input
rlabel metal3 s 100 140112 400 140168 6 state[59]
port 340 nsew signal input
rlabel metal3 s 249600 7056 249900 7112 6 state[5]
port 341 nsew signal input
rlabel metal2 s 38640 100 38696 400 6 state[60]
port 342 nsew signal input
rlabel metal2 s 121968 100 122024 400 6 state[61]
port 343 nsew signal input
rlabel metal3 s 249600 105504 249900 105560 6 state[62]
port 344 nsew signal input
rlabel metal2 s 201600 249600 201656 249900 6 state[63]
port 345 nsew signal input
rlabel metal3 s 249600 220080 249900 220136 6 state[64]
port 346 nsew signal input
rlabel metal3 s 249600 12096 249900 12152 6 state[65]
port 347 nsew signal input
rlabel metal2 s 20496 100 20552 400 6 state[66]
port 348 nsew signal input
rlabel metal3 s 249600 139440 249900 139496 6 state[67]
port 349 nsew signal input
rlabel metal2 s 5040 100 5096 400 6 state[68]
port 350 nsew signal input
rlabel metal3 s 249600 227808 249900 227864 6 state[69]
port 351 nsew signal input
rlabel metal2 s 191520 249600 191576 249900 6 state[6]
port 352 nsew signal input
rlabel metal3 s 249600 27888 249900 27944 6 state[70]
port 353 nsew signal input
rlabel metal2 s 183456 249600 183512 249900 6 state[71]
port 354 nsew signal input
rlabel metal2 s 168672 100 168728 400 6 state[72]
port 355 nsew signal input
rlabel metal3 s 100 82992 400 83048 6 state[73]
port 356 nsew signal input
rlabel metal2 s 165984 100 166040 400 6 state[74]
port 357 nsew signal input
rlabel metal2 s 0 100 56 400 6 state[75]
port 358 nsew signal input
rlabel metal2 s 197232 100 197288 400 6 state[76]
port 359 nsew signal input
rlabel metal3 s 100 124656 400 124712 6 state[77]
port 360 nsew signal input
rlabel metal3 s 100 220752 400 220808 6 state[78]
port 361 nsew signal input
rlabel metal2 s 71904 249600 71960 249900 6 state[79]
port 362 nsew signal input
rlabel metal3 s 100 85680 400 85736 6 state[7]
port 363 nsew signal input
rlabel metal2 s 51744 100 51800 400 6 state[80]
port 364 nsew signal input
rlabel metal2 s 18144 100 18200 400 6 state[81]
port 365 nsew signal input
rlabel metal2 s 131712 249600 131768 249900 6 state[82]
port 366 nsew signal input
rlabel metal2 s 76944 249600 77000 249900 6 state[83]
port 367 nsew signal input
rlabel metal2 s 134736 100 134792 400 6 state[84]
port 368 nsew signal input
rlabel metal2 s 175728 249600 175784 249900 6 state[85]
port 369 nsew signal input
rlabel metal3 s 249600 69216 249900 69272 6 state[86]
port 370 nsew signal input
rlabel metal3 s 100 165984 400 166040 6 state[87]
port 371 nsew signal input
rlabel metal3 s 249600 191520 249900 191576 6 state[88]
port 372 nsew signal input
rlabel metal2 s 54432 100 54488 400 6 state[89]
port 373 nsew signal input
rlabel metal2 s 96096 100 96152 400 6 state[8]
port 374 nsew signal input
rlabel metal3 s 100 23184 400 23240 6 state[90]
port 375 nsew signal input
rlabel metal3 s 249600 183456 249900 183512 6 state[91]
port 376 nsew signal input
rlabel metal2 s 150528 100 150584 400 6 state[92]
port 377 nsew signal input
rlabel metal2 s 165312 249600 165368 249900 6 state[93]
port 378 nsew signal input
rlabel metal2 s 162960 249600 163016 249900 6 state[94]
port 379 nsew signal input
rlabel metal3 s 100 230832 400 230888 6 state[95]
port 380 nsew signal input
rlabel metal2 s 27888 249600 27944 249900 6 state[96]
port 381 nsew signal input
rlabel metal2 s 181776 100 181832 400 6 state[97]
port 382 nsew signal input
rlabel metal3 s 100 54432 400 54488 6 state[98]
port 383 nsew signal input
rlabel metal3 s 100 207648 400 207704 6 state[99]
port 384 nsew signal input
rlabel metal3 s 249600 123984 249900 124040 6 state[9]
port 385 nsew signal input
rlabel metal4 s 2224 1538 2384 248166 6 vdd
port 386 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 248166 6 vdd
port 386 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 248166 6 vdd
port 386 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 248166 6 vdd
port 386 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 248166 6 vdd
port 386 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 248166 6 vdd
port 386 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 248166 6 vdd
port 386 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 248166 6 vdd
port 386 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 248166 6 vdd
port 386 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 248166 6 vdd
port 386 nsew power bidirectional
rlabel metal4 s 155824 1538 155984 248166 6 vdd
port 386 nsew power bidirectional
rlabel metal4 s 171184 1538 171344 248166 6 vdd
port 386 nsew power bidirectional
rlabel metal4 s 186544 1538 186704 248166 6 vdd
port 386 nsew power bidirectional
rlabel metal4 s 201904 1538 202064 248166 6 vdd
port 386 nsew power bidirectional
rlabel metal4 s 217264 1538 217424 248166 6 vdd
port 386 nsew power bidirectional
rlabel metal4 s 232624 1538 232784 248166 6 vdd
port 386 nsew power bidirectional
rlabel metal4 s 247984 1538 248144 248166 6 vdd
port 386 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 248166 6 vss
port 387 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 248166 6 vss
port 387 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 248166 6 vss
port 387 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 248166 6 vss
port 387 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 248166 6 vss
port 387 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 248166 6 vss
port 387 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 248166 6 vss
port 387 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 248166 6 vss
port 387 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 248166 6 vss
port 387 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 248166 6 vss
port 387 nsew ground bidirectional
rlabel metal4 s 163504 1538 163664 248166 6 vss
port 387 nsew ground bidirectional
rlabel metal4 s 178864 1538 179024 248166 6 vss
port 387 nsew ground bidirectional
rlabel metal4 s 194224 1538 194384 248166 6 vss
port 387 nsew ground bidirectional
rlabel metal4 s 209584 1538 209744 248166 6 vss
port 387 nsew ground bidirectional
rlabel metal4 s 224944 1538 225104 248166 6 vss
port 387 nsew ground bidirectional
rlabel metal4 s 240304 1538 240464 248166 6 vss
port 387 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 250000 250000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 94083646
string GDS_FILE /home/urielcho/Proyectos_caravel/gf180nm/aes128/openlane/aes128/runs/22_12_05_01_35/results/signoff/aes128.magic.gds
string GDS_START 326160
<< end >>

