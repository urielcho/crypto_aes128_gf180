VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO aes128
  CLASS BLOCK ;
  FOREIGN aes128 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2500.000 BY 2500.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1038.240 4.000 1038.800 ;
    END
  END clk
  PIN key[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2328.480 2496.000 2329.040 2499.000 ;
    END
  END key[0]
  PIN key[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 594.720 4.000 595.280 ;
    END
  END key[100]
  PIN key[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2042.880 2496.000 2043.440 2499.000 ;
    END
  END key[101]
  PIN key[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 154.560 4.000 155.120 ;
    END
  END key[102]
  PIN key[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1505.280 4.000 1505.840 ;
    END
  END key[103]
  PIN key[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1374.240 4.000 1374.800 ;
    END
  END key[104]
  PIN key[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 460.320 2499.000 460.880 ;
    END
  END key[105]
  PIN key[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 2180.640 4.000 2181.200 ;
    END
  END key[106]
  PIN key[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1004.640 2496.000 1005.200 2499.000 ;
    END
  END key[107]
  PIN key[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 850.080 2496.000 850.640 2499.000 ;
    END
  END key[108]
  PIN key[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1706.880 2496.000 1707.440 2499.000 ;
    END
  END key[109]
  PIN key[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 564.480 2499.000 565.040 ;
    END
  END key[10]
  PIN key[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2224.320 2496.000 2224.880 2499.000 ;
    END
  END key[110]
  PIN key[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1609.440 4.000 1610.000 ;
    END
  END key[111]
  PIN key[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1323.840 1.000 1324.400 4.000 ;
    END
  END key[112]
  PIN key[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 796.320 2499.000 796.880 ;
    END
  END key[113]
  PIN key[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2405.760 2496.000 2406.320 2499.000 ;
    END
  END key[114]
  PIN key[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1999.200 4.000 1999.760 ;
    END
  END key[115]
  PIN key[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 648.480 4.000 649.040 ;
    END
  END key[116]
  PIN key[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2355.360 2499.000 2355.920 ;
    END
  END key[117]
  PIN key[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1498.560 2499.000 1499.120 ;
    END
  END key[118]
  PIN key[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2257.920 1.000 2258.480 4.000 ;
    END
  END key[119]
  PIN key[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1938.720 2496.000 1939.280 2499.000 ;
    END
  END key[11]
  PIN key[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1582.560 1.000 1583.120 4.000 ;
    END
  END key[120]
  PIN key[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 2439.360 4.000 2439.920 ;
    END
  END key[121]
  PIN key[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 954.240 2496.000 954.800 2499.000 ;
    END
  END key[122]
  PIN key[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2120.160 2499.000 2120.720 ;
    END
  END key[123]
  PIN key[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 900.480 2499.000 901.040 ;
    END
  END key[124]
  PIN key[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 2388.960 4.000 2389.520 ;
    END
  END key[125]
  PIN key[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1861.440 2496.000 1862.000 2499.000 ;
    END
  END key[126]
  PIN key[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1811.040 2499.000 1811.600 ;
    END
  END key[127]
  PIN key[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 571.200 1.000 571.760 4.000 ;
    END
  END key[12]
  PIN key[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1317.120 2499.000 1317.680 ;
    END
  END key[13]
  PIN key[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 1.000 155.120 4.000 ;
    END
  END key[14]
  PIN key[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2439.360 1.000 2439.920 4.000 ;
    END
  END key[15]
  PIN key[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1532.160 1.000 1532.720 4.000 ;
    END
  END key[16]
  PIN key[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 776.160 4.000 776.720 ;
    END
  END key[17]
  PIN key[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 803.040 4.000 803.600 ;
    END
  END key[18]
  PIN key[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 588.000 2499.000 588.560 ;
    END
  END key[19]
  PIN key[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2328.480 2499.000 2329.040 ;
    END
  END key[1]
  PIN key[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2207.520 1.000 2208.080 4.000 ;
    END
  END key[20]
  PIN key[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1680.000 2499.000 1680.560 ;
    END
  END key[21]
  PIN key[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2486.400 2499.000 2486.960 ;
    END
  END key[22]
  PIN key[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1632.960 1.000 1633.520 4.000 ;
    END
  END key[23]
  PIN key[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 204.960 4.000 205.520 ;
    END
  END key[24]
  PIN key[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 614.880 2496.000 615.440 2499.000 ;
    END
  END key[25]
  PIN key[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 564.480 2496.000 565.040 2499.000 ;
    END
  END key[26]
  PIN key[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1263.360 2496.000 1263.920 2499.000 ;
    END
  END key[27]
  PIN key[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1868.160 4.000 1868.720 ;
    END
  END key[28]
  PIN key[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 231.840 1.000 232.400 4.000 ;
    END
  END key[29]
  PIN key[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1992.480 2499.000 1993.040 ;
    END
  END key[2]
  PIN key[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1212.960 2499.000 1213.520 ;
    END
  END key[30]
  PIN key[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 2496.000 94.640 2499.000 ;
    END
  END key[31]
  PIN key[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2335.200 1.000 2335.760 4.000 ;
    END
  END key[32]
  PIN key[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 329.280 2499.000 329.840 ;
    END
  END key[33]
  PIN key[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1548.960 2499.000 1549.520 ;
    END
  END key[34]
  PIN key[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 386.400 4.000 386.960 ;
    END
  END key[35]
  PIN key[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2459.520 2499.000 2460.080 ;
    END
  END key[36]
  PIN key[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1108.800 2499.000 1109.360 ;
    END
  END key[37]
  PIN key[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2224.320 2499.000 2224.880 ;
    END
  END key[38]
  PIN key[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1817.760 4.000 1818.320 ;
    END
  END key[39]
  PIN key[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1602.720 2496.000 1603.280 2499.000 ;
    END
  END key[3]
  PIN key[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1945.440 4.000 1946.000 ;
    END
  END key[40]
  PIN key[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 594.720 1.000 595.280 4.000 ;
    END
  END key[41]
  PIN key[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2153.760 1.000 2154.320 4.000 ;
    END
  END key[42]
  PIN key[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1212.960 2496.000 1213.520 2499.000 ;
    END
  END key[43]
  PIN key[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1764.000 1.000 1764.560 4.000 ;
    END
  END key[44]
  PIN key[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1992.480 2496.000 1993.040 2499.000 ;
    END
  END key[45]
  PIN key[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2412.480 1.000 2413.040 4.000 ;
    END
  END key[46]
  PIN key[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1401.120 1.000 1401.680 4.000 ;
    END
  END key[47]
  PIN key[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1444.800 2496.000 1445.360 2499.000 ;
    END
  END key[48]
  PIN key[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1270.080 1.000 1270.640 4.000 ;
    END
  END key[49]
  PIN key[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2016.000 2499.000 2016.560 ;
    END
  END key[4]
  PIN key[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1055.040 2496.000 1055.600 2499.000 ;
    END
  END key[50]
  PIN key[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1290.240 2499.000 1290.800 ;
    END
  END key[51]
  PIN key[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1945.440 1.000 1946.000 4.000 ;
    END
  END key[52]
  PIN key[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1888.320 2499.000 1888.880 ;
    END
  END key[53]
  PIN key[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1861.440 2499.000 1862.000 ;
    END
  END key[54]
  PIN key[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1088.640 1.000 1089.200 4.000 ;
    END
  END key[55]
  PIN key[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 285.600 1.000 286.160 4.000 ;
    END
  END key[56]
  PIN key[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1632.960 4.000 1633.520 ;
    END
  END key[57]
  PIN key[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 483.840 2499.000 484.400 ;
    END
  END key[58]
  PIN key[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 483.840 2496.000 484.400 2499.000 ;
    END
  END key[59]
  PIN key[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1999.200 1.000 1999.760 4.000 ;
    END
  END key[5]
  PIN key[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 43.680 2499.000 44.240 ;
    END
  END key[60]
  PIN key[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 2496.000 44.240 2499.000 ;
    END
  END key[61]
  PIN key[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 934.080 4.000 934.640 ;
    END
  END key[62]
  PIN key[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2382.240 2499.000 2382.800 ;
    END
  END key[63]
  PIN key[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 934.080 1.000 934.640 4.000 ;
    END
  END key[64]
  PIN key[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1165.920 1.000 1166.480 4.000 ;
    END
  END key[65]
  PIN key[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 406.560 2496.000 407.120 2499.000 ;
    END
  END key[66]
  PIN key[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2173.920 2499.000 2174.480 ;
    END
  END key[67]
  PIN key[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 641.760 2496.000 642.320 2499.000 ;
    END
  END key[68]
  PIN key[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 2496.000 148.400 2499.000 ;
    END
  END key[69]
  PIN key[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1895.040 4.000 1895.600 ;
    END
  END key[6]
  PIN key[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 356.160 2496.000 356.720 2499.000 ;
    END
  END key[70]
  PIN key[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 614.880 2499.000 615.440 ;
    END
  END key[71]
  PIN key[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 752.640 1.000 753.200 4.000 ;
    END
  END key[72]
  PIN key[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1135.680 2496.000 1136.240 2499.000 ;
    END
  END key[73]
  PIN key[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 621.600 4.000 622.160 ;
    END
  END key[74]
  PIN key[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1239.840 2496.000 1240.400 2499.000 ;
    END
  END key[75]
  PIN key[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 252.000 2499.000 252.560 ;
    END
  END key[76]
  PIN key[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 648.480 1.000 649.040 4.000 ;
    END
  END key[77]
  PIN key[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1471.680 2496.000 1472.240 2499.000 ;
    END
  END key[78]
  PIN key[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1706.880 2499.000 1707.440 ;
    END
  END key[79]
  PIN key[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 174.720 2499.000 175.280 ;
    END
  END key[7]
  PIN key[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2486.400 2496.000 2486.960 2499.000 ;
    END
  END key[80]
  PIN key[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1428.000 4.000 1428.560 ;
    END
  END key[81]
  PIN key[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1498.560 2496.000 1499.120 2499.000 ;
    END
  END key[82]
  PIN key[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2173.920 2496.000 2174.480 2499.000 ;
    END
  END key[83]
  PIN key[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2069.760 2499.000 2070.320 ;
    END
  END key[84]
  PIN key[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 285.600 4.000 286.160 ;
    END
  END key[85]
  PIN key[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2042.880 2499.000 2043.440 ;
    END
  END key[86]
  PIN key[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1088.640 4.000 1089.200 ;
    END
  END key[87]
  PIN key[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 490.560 1.000 491.120 4.000 ;
    END
  END key[88]
  PIN key[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 252.000 2496.000 252.560 2499.000 ;
    END
  END key[89]
  PIN key[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1737.120 4.000 1737.680 ;
    END
  END key[8]
  PIN key[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1038.240 1.000 1038.800 4.000 ;
    END
  END key[90]
  PIN key[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 829.920 1.000 830.480 4.000 ;
    END
  END key[91]
  PIN key[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 362.880 1.000 363.440 4.000 ;
    END
  END key[92]
  PIN key[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2180.640 1.000 2181.200 4.000 ;
    END
  END key[93]
  PIN key[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 698.880 1.000 699.440 4.000 ;
    END
  END key[94]
  PIN key[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 2493.120 4.000 2493.680 ;
    END
  END key[95]
  PIN key[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1764.000 4.000 1764.560 ;
    END
  END key[96]
  PIN key[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 745.920 2496.000 746.480 2499.000 ;
    END
  END key[97]
  PIN key[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 752.640 4.000 753.200 ;
    END
  END key[98]
  PIN key[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1159.200 2496.000 1159.760 2499.000 ;
    END
  END key[99]
  PIN key[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 954.240 2499.000 954.800 ;
    END
  END key[9]
  PIN out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1011.360 1.000 1011.920 4.000 ;
    END
  END out[0]
  PIN out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 406.560 2499.000 407.120 ;
    END
  END out[100]
  PIN out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 2496.000 17.360 2499.000 ;
    END
  END out[101]
  PIN out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 302.400 2499.000 302.960 ;
    END
  END out[102]
  PIN out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 725.760 4.000 726.320 ;
    END
  END out[103]
  PIN out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 50.400 4.000 50.960 ;
    END
  END out[104]
  PIN out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2284.800 1.000 2285.360 4.000 ;
    END
  END out[105]
  PIN out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 803.040 1.000 803.600 4.000 ;
    END
  END out[106]
  PIN out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2096.640 2496.000 2097.200 2499.000 ;
    END
  END out[107]
  PIN out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1532.160 4.000 1532.720 ;
    END
  END out[108]
  PIN out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 198.240 2496.000 198.800 2499.000 ;
    END
  END out[109]
  PIN out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1142.400 1.000 1142.960 4.000 ;
    END
  END out[10]
  PIN out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 2362.080 4.000 2362.640 ;
    END
  END out[110]
  PIN out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1394.400 2496.000 1394.960 2499.000 ;
    END
  END out[111]
  PIN out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1525.440 2496.000 1526.000 2499.000 ;
    END
  END out[112]
  PIN out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 537.600 2499.000 538.160 ;
    END
  END out[113]
  PIN out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2251.200 2499.000 2251.760 ;
    END
  END out[114]
  PIN out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2049.600 1.000 2050.160 4.000 ;
    END
  END out[115]
  PIN out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 873.600 2499.000 874.160 ;
    END
  END out[116]
  PIN out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 927.360 2499.000 927.920 ;
    END
  END out[117]
  PIN out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1609.440 1.000 1610.000 4.000 ;
    END
  END out[118]
  PIN out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 725.760 1.000 726.320 4.000 ;
    END
  END out[119]
  PIN out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 856.800 1.000 857.360 4.000 ;
    END
  END out[11]
  PIN out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 668.640 2499.000 669.200 ;
    END
  END out[120]
  PIN out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1965.600 2499.000 1966.160 ;
    END
  END out[121]
  PIN out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1790.880 4.000 1791.440 ;
    END
  END out[122]
  PIN out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 413.280 1.000 413.840 4.000 ;
    END
  END out[123]
  PIN out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1629.600 2499.000 1630.160 ;
    END
  END out[124]
  PIN out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1555.680 4.000 1556.240 ;
    END
  END out[125]
  PIN out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 823.200 2499.000 823.760 ;
    END
  END out[126]
  PIN out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 120.960 2496.000 121.520 2499.000 ;
    END
  END out[127]
  PIN out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1367.520 2499.000 1368.080 ;
    END
  END out[12]
  PIN out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1548.960 2496.000 1549.520 2499.000 ;
    END
  END out[13]
  PIN out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 181.440 4.000 182.000 ;
    END
  END out[14]
  PIN out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 433.440 2499.000 434.000 ;
    END
  END out[15]
  PIN out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1344.000 2496.000 1344.560 2499.000 ;
    END
  END out[16]
  PIN out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 440.160 4.000 440.720 ;
    END
  END out[17]
  PIN out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 537.600 2496.000 538.160 2499.000 ;
    END
  END out[18]
  PIN out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1602.720 2499.000 1603.280 ;
    END
  END out[19]
  PIN out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 984.480 1.000 985.040 4.000 ;
    END
  END out[1]
  PIN out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 880.320 1.000 880.880 4.000 ;
    END
  END out[20]
  PIN out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 850.080 2499.000 850.640 ;
    END
  END out[21]
  PIN out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 796.320 2496.000 796.880 2499.000 ;
    END
  END out[22]
  PIN out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 383.040 2496.000 383.600 2499.000 ;
    END
  END out[23]
  PIN out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 225.120 2499.000 225.680 ;
    END
  END out[24]
  PIN out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1115.520 1.000 1116.080 4.000 ;
    END
  END out[25]
  PIN out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2200.800 2496.000 2201.360 2499.000 ;
    END
  END out[26]
  PIN out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1653.120 2499.000 1653.680 ;
    END
  END out[27]
  PIN out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 413.280 4.000 413.840 ;
    END
  END out[28]
  PIN out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 2412.480 4.000 2413.040 ;
    END
  END out[29]
  PIN out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1011.360 4.000 1011.920 ;
    END
  END out[2]
  PIN out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1451.520 1.000 1452.080 4.000 ;
    END
  END out[30]
  PIN out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 588.000 2496.000 588.560 2499.000 ;
    END
  END out[31]
  PIN out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2120.160 2496.000 2120.720 2499.000 ;
    END
  END out[32]
  PIN out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1757.280 2499.000 1757.840 ;
    END
  END out[33]
  PIN out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 1.000 128.240 4.000 ;
    END
  END out[34]
  PIN out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 2103.360 4.000 2103.920 ;
    END
  END out[35]
  PIN out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 174.720 2496.000 175.280 2499.000 ;
    END
  END out[36]
  PIN out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1575.840 2496.000 1576.400 2499.000 ;
    END
  END out[37]
  PIN out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1921.920 4.000 1922.480 ;
    END
  END out[38]
  PIN out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 336.000 4.000 336.560 ;
    END
  END out[39]
  PIN out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2103.360 1.000 2103.920 4.000 ;
    END
  END out[3]
  PIN out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1031.520 2499.000 1032.080 ;
    END
  END out[40]
  PIN out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 94.080 2499.000 94.640 ;
    END
  END out[41]
  PIN out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 77.280 4.000 77.840 ;
    END
  END out[42]
  PIN out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1108.800 2496.000 1109.360 2499.000 ;
    END
  END out[43]
  PIN out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1296.960 1.000 1297.520 4.000 ;
    END
  END out[44]
  PIN out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 2466.240 4.000 2466.800 ;
    END
  END out[45]
  PIN out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1192.800 1.000 1193.360 4.000 ;
    END
  END out[46]
  PIN out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 383.040 2499.000 383.600 ;
    END
  END out[47]
  PIN out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2251.200 2496.000 2251.760 2499.000 ;
    END
  END out[48]
  PIN out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 490.560 4.000 491.120 ;
    END
  END out[49]
  PIN out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1421.280 2496.000 1421.840 2499.000 ;
    END
  END out[4]
  PIN out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 880.320 4.000 880.880 ;
    END
  END out[50]
  PIN out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2355.360 2496.000 2355.920 2499.000 ;
    END
  END out[51]
  PIN out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 433.440 2496.000 434.000 2499.000 ;
    END
  END out[52]
  PIN out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 672.000 4.000 672.560 ;
    END
  END out[53]
  PIN out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 16.800 2499.000 17.360 ;
    END
  END out[54]
  PIN out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 2284.800 4.000 2285.360 ;
    END
  END out[55]
  PIN out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 2126.880 4.000 2127.440 ;
    END
  END out[56]
  PIN out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1478.400 1.000 1478.960 4.000 ;
    END
  END out[57]
  PIN out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 977.760 2499.000 978.320 ;
    END
  END out[58]
  PIN out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 745.920 2499.000 746.480 ;
    END
  END out[59]
  PIN out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 873.600 2496.000 874.160 2499.000 ;
    END
  END out[5]
  PIN out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1186.080 2499.000 1186.640 ;
    END
  END out[60]
  PIN out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1790.880 1.000 1791.440 4.000 ;
    END
  END out[61]
  PIN out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 23.520 4.000 24.080 ;
    END
  END out[62]
  PIN out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1737.120 1.000 1737.680 4.000 ;
    END
  END out[63]
  PIN out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2076.480 1.000 2077.040 4.000 ;
    END
  END out[64]
  PIN out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 336.000 1.000 336.560 4.000 ;
    END
  END out[65]
  PIN out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1686.720 4.000 1687.280 ;
    END
  END out[66]
  PIN out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1895.040 1.000 1895.600 4.000 ;
    END
  END out[67]
  PIN out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1165.920 4.000 1166.480 ;
    END
  END out[68]
  PIN out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1841.280 4.000 1841.840 ;
    END
  END out[69]
  PIN out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2432.640 2499.000 2433.200 ;
    END
  END out[6]
  PIN out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 517.440 4.000 518.000 ;
    END
  END out[70]
  PIN out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1347.360 4.000 1347.920 ;
    END
  END out[71]
  PIN out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 672.000 1.000 672.560 4.000 ;
    END
  END out[72]
  PIN out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1344.000 2499.000 1344.560 ;
    END
  END out[73]
  PIN out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2126.880 1.000 2127.440 4.000 ;
    END
  END out[74]
  PIN out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1965.600 2496.000 1966.160 2499.000 ;
    END
  END out[75]
  PIN out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 440.160 1.000 440.720 4.000 ;
    END
  END out[76]
  PIN out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 510.720 2496.000 511.280 2499.000 ;
    END
  END out[77]
  PIN out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2147.040 2499.000 2147.600 ;
    END
  END out[78]
  PIN out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 907.200 4.000 907.760 ;
    END
  END out[79]
  PIN out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1938.720 2499.000 1939.280 ;
    END
  END out[7]
  PIN out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1367.520 2496.000 1368.080 2499.000 ;
    END
  END out[80]
  PIN out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 258.720 4.000 259.280 ;
    END
  END out[81]
  PIN out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1115.520 4.000 1116.080 ;
    END
  END out[82]
  PIN out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1478.400 4.000 1478.960 ;
    END
  END out[83]
  PIN out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1081.920 2496.000 1082.480 2499.000 ;
    END
  END out[84]
  PIN out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 1.000 24.080 4.000 ;
    END
  END out[85]
  PIN out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 692.160 2496.000 692.720 2499.000 ;
    END
  END out[86]
  PIN out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1246.560 1.000 1247.120 4.000 ;
    END
  END out[87]
  PIN out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2493.120 1.000 2493.680 4.000 ;
    END
  END out[88]
  PIN out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2405.760 2499.000 2406.320 ;
    END
  END out[89]
  PIN out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 198.240 2499.000 198.800 ;
    END
  END out[8]
  PIN out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1186.080 2496.000 1186.640 2499.000 ;
    END
  END out[90]
  PIN out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 1.000 77.840 4.000 ;
    END
  END out[91]
  PIN out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 467.040 1.000 467.600 4.000 ;
    END
  END out[92]
  PIN out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1061.760 1.000 1062.320 4.000 ;
    END
  END out[93]
  PIN out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2278.080 2496.000 2278.640 2499.000 ;
    END
  END out[94]
  PIN out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 2022.720 4.000 2023.280 ;
    END
  END out[95]
  PIN out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 907.200 1.000 907.760 4.000 ;
    END
  END out[96]
  PIN out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 100.800 4.000 101.360 ;
    END
  END out[97]
  PIN out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1081.920 2499.000 1082.480 ;
    END
  END out[98]
  PIN out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 2257.920 4.000 2258.480 ;
    END
  END out[99]
  PIN out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1868.160 1.000 1868.720 4.000 ;
    END
  END out[9]
  PIN state[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 127.680 4.000 128.240 ;
    END
  END state[0]
  PIN state[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2388.960 1.000 2389.520 4.000 ;
    END
  END state[100]
  PIN state[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1444.800 2499.000 1445.360 ;
    END
  END state[101]
  PIN state[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1888.320 2496.000 1888.880 2499.000 ;
    END
  END state[102]
  PIN state[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1159.200 2499.000 1159.760 ;
    END
  END state[103]
  PIN state[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1972.320 4.000 1972.880 ;
    END
  END state[104]
  PIN state[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1451.520 4.000 1452.080 ;
    END
  END state[105]
  PIN state[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 147.840 2499.000 148.400 ;
    END
  END state[106]
  PIN state[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1680.000 2496.000 1680.560 2499.000 ;
    END
  END state[107]
  PIN state[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2231.040 1.000 2231.600 4.000 ;
    END
  END state[108]
  PIN state[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 302.400 2496.000 302.960 2499.000 ;
    END
  END state[109]
  PIN state[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 309.120 1.000 309.680 4.000 ;
    END
  END state[10]
  PIN state[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1135.680 2499.000 1136.240 ;
    END
  END state[110]
  PIN state[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 2496.000 71.120 2499.000 ;
    END
  END state[111]
  PIN state[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1525.440 2499.000 1526.000 ;
    END
  END state[112]
  PIN state[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 621.600 1.000 622.160 4.000 ;
    END
  END state[113]
  PIN state[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2308.320 1.000 2308.880 4.000 ;
    END
  END state[114]
  PIN state[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 927.360 2496.000 927.920 2499.000 ;
    END
  END state[115]
  PIN state[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2304.960 2496.000 2305.520 2499.000 ;
    END
  END state[116]
  PIN state[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1784.160 2499.000 1784.720 ;
    END
  END state[117]
  PIN state[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 823.200 2496.000 823.760 2499.000 ;
    END
  END state[118]
  PIN state[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1031.520 2496.000 1032.080 2499.000 ;
    END
  END state[119]
  PIN state[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 356.160 2499.000 356.720 ;
    END
  END state[11]
  PIN state[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1323.840 4.000 1324.400 ;
    END
  END state[120]
  PIN state[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1192.800 4.000 1193.360 ;
    END
  END state[121]
  PIN state[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1811.040 2496.000 1811.600 2499.000 ;
    END
  END state[122]
  PIN state[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1290.240 2496.000 1290.800 2499.000 ;
    END
  END state[123]
  PIN state[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 329.280 2496.000 329.840 2499.000 ;
    END
  END state[124]
  PIN state[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 984.480 4.000 985.040 ;
    END
  END state[125]
  PIN state[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 2335.200 4.000 2335.760 ;
    END
  END state[126]
  PIN state[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1730.400 2499.000 1730.960 ;
    END
  END state[127]
  PIN state[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1575.840 2499.000 1576.400 ;
    END
  END state[12]
  PIN state[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1555.680 1.000 1556.240 4.000 ;
    END
  END state[13]
  PIN state[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1421.280 2499.000 1421.840 ;
    END
  END state[14]
  PIN state[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1219.680 4.000 1220.240 ;
    END
  END state[15]
  PIN state[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2362.080 1.000 2362.640 4.000 ;
    END
  END state[16]
  PIN state[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1730.400 2496.000 1730.960 2499.000 ;
    END
  END state[17]
  PIN state[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2432.640 2496.000 2433.200 2499.000 ;
    END
  END state[18]
  PIN state[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1374.240 1.000 1374.800 4.000 ;
    END
  END state[19]
  PIN state[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 698.880 4.000 699.440 ;
    END
  END state[1]
  PIN state[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 510.720 2499.000 511.280 ;
    END
  END state[20]
  PIN state[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 460.320 2496.000 460.880 2499.000 ;
    END
  END state[21]
  PIN state[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 467.040 4.000 467.600 ;
    END
  END state[22]
  PIN state[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 258.720 1.000 259.280 4.000 ;
    END
  END state[23]
  PIN state[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 977.760 2496.000 978.320 2499.000 ;
    END
  END state[24]
  PIN state[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 960.960 4.000 961.520 ;
    END
  END state[25]
  PIN state[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2304.960 2499.000 2305.520 ;
    END
  END state[26]
  PIN state[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 309.120 4.000 309.680 ;
    END
  END state[27]
  PIN state[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2069.760 2496.000 2070.320 2499.000 ;
    END
  END state[28]
  PIN state[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1004.640 2499.000 1005.200 ;
    END
  END state[29]
  PIN state[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1921.920 1.000 1922.480 4.000 ;
    END
  END state[2]
  PIN state[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1061.760 4.000 1062.320 ;
    END
  END state[30]
  PIN state[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1841.280 1.000 1841.840 4.000 ;
    END
  END state[31]
  PIN state[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1296.960 4.000 1297.520 ;
    END
  END state[32]
  PIN state[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1713.600 4.000 1714.160 ;
    END
  END state[33]
  PIN state[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2466.240 1.000 2466.800 4.000 ;
    END
  END state[34]
  PIN state[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 641.760 2499.000 642.320 ;
    END
  END state[35]
  PIN state[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 900.480 2496.000 901.040 2499.000 ;
    END
  END state[36]
  PIN state[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2096.640 2499.000 2097.200 ;
    END
  END state[37]
  PIN state[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 2049.600 4.000 2050.160 ;
    END
  END state[38]
  PIN state[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 2231.040 4.000 2231.600 ;
    END
  END state[39]
  PIN state[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 2153.760 4.000 2154.320 ;
    END
  END state[3]
  PIN state[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 1.000 101.360 4.000 ;
    END
  END state[40]
  PIN state[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 571.200 4.000 571.760 ;
    END
  END state[41]
  PIN state[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1263.360 2499.000 1263.920 ;
    END
  END state[42]
  PIN state[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1428.000 1.000 1428.560 4.000 ;
    END
  END state[43]
  PIN state[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1784.160 2496.000 1784.720 2499.000 ;
    END
  END state[44]
  PIN state[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2382.240 2496.000 2382.800 2499.000 ;
    END
  END state[45]
  PIN state[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 225.120 2496.000 225.680 2499.000 ;
    END
  END state[46]
  PIN state[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1142.400 4.000 1142.960 ;
    END
  END state[47]
  PIN state[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1270.080 4.000 1270.640 ;
    END
  END state[48]
  PIN state[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2459.520 2496.000 2460.080 2499.000 ;
    END
  END state[49]
  PIN state[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1582.560 4.000 1583.120 ;
    END
  END state[4]
  PIN state[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 362.880 4.000 363.440 ;
    END
  END state[50]
  PIN state[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 769.440 2499.000 770.000 ;
    END
  END state[51]
  PIN state[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1713.600 1.000 1714.160 4.000 ;
    END
  END state[52]
  PIN state[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2147.040 2496.000 2147.600 2499.000 ;
    END
  END state[53]
  PIN state[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 668.640 2496.000 669.200 2499.000 ;
    END
  END state[54]
  PIN state[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 776.160 1.000 776.720 4.000 ;
    END
  END state[55]
  PIN state[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1471.680 2499.000 1472.240 ;
    END
  END state[56]
  PIN state[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2022.720 1.000 2023.280 4.000 ;
    END
  END state[57]
  PIN state[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 719.040 2499.000 719.600 ;
    END
  END state[58]
  PIN state[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1401.120 4.000 1401.680 ;
    END
  END state[59]
  PIN state[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 70.560 2499.000 71.120 ;
    END
  END state[5]
  PIN state[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 386.400 1.000 386.960 4.000 ;
    END
  END state[60]
  PIN state[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1219.680 1.000 1220.240 4.000 ;
    END
  END state[61]
  PIN state[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1055.040 2499.000 1055.600 ;
    END
  END state[62]
  PIN state[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2016.000 2496.000 2016.560 2499.000 ;
    END
  END state[63]
  PIN state[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2200.800 2499.000 2201.360 ;
    END
  END state[64]
  PIN state[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 120.960 2499.000 121.520 ;
    END
  END state[65]
  PIN state[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 1.000 205.520 4.000 ;
    END
  END state[66]
  PIN state[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1394.400 2499.000 1394.960 ;
    END
  END state[67]
  PIN state[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 1.000 50.960 4.000 ;
    END
  END state[68]
  PIN state[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2278.080 2499.000 2278.640 ;
    END
  END state[69]
  PIN state[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1915.200 2496.000 1915.760 2499.000 ;
    END
  END state[6]
  PIN state[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 278.880 2499.000 279.440 ;
    END
  END state[70]
  PIN state[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1834.560 2496.000 1835.120 2499.000 ;
    END
  END state[71]
  PIN state[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1686.720 1.000 1687.280 4.000 ;
    END
  END state[72]
  PIN state[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 829.920 4.000 830.480 ;
    END
  END state[73]
  PIN state[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1659.840 1.000 1660.400 4.000 ;
    END
  END state[74]
  PIN state[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1.000 0.560 4.000 ;
    END
  END state[75]
  PIN state[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1972.320 1.000 1972.880 4.000 ;
    END
  END state[76]
  PIN state[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1246.560 4.000 1247.120 ;
    END
  END state[77]
  PIN state[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 2207.520 4.000 2208.080 ;
    END
  END state[78]
  PIN state[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 719.040 2496.000 719.600 2499.000 ;
    END
  END state[79]
  PIN state[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 856.800 4.000 857.360 ;
    END
  END state[7]
  PIN state[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 517.440 1.000 518.000 4.000 ;
    END
  END state[80]
  PIN state[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 181.440 1.000 182.000 4.000 ;
    END
  END state[81]
  PIN state[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1317.120 2496.000 1317.680 2499.000 ;
    END
  END state[82]
  PIN state[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 769.440 2496.000 770.000 2499.000 ;
    END
  END state[83]
  PIN state[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1347.360 1.000 1347.920 4.000 ;
    END
  END state[84]
  PIN state[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1757.280 2496.000 1757.840 2499.000 ;
    END
  END state[85]
  PIN state[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 692.160 2499.000 692.720 ;
    END
  END state[86]
  PIN state[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1659.840 4.000 1660.400 ;
    END
  END state[87]
  PIN state[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1915.200 2499.000 1915.760 ;
    END
  END state[88]
  PIN state[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 544.320 1.000 544.880 4.000 ;
    END
  END state[89]
  PIN state[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 960.960 1.000 961.520 4.000 ;
    END
  END state[8]
  PIN state[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 231.840 4.000 232.400 ;
    END
  END state[90]
  PIN state[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1834.560 2499.000 1835.120 ;
    END
  END state[91]
  PIN state[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1505.280 1.000 1505.840 4.000 ;
    END
  END state[92]
  PIN state[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1653.120 2496.000 1653.680 2499.000 ;
    END
  END state[93]
  PIN state[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1629.600 2496.000 1630.160 2499.000 ;
    END
  END state[94]
  PIN state[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 2308.320 4.000 2308.880 ;
    END
  END state[95]
  PIN state[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 278.880 2496.000 279.440 2499.000 ;
    END
  END state[96]
  PIN state[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1817.760 1.000 1818.320 4.000 ;
    END
  END state[97]
  PIN state[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 544.320 4.000 544.880 ;
    END
  END state[98]
  PIN state[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 2076.480 4.000 2077.040 ;
    END
  END state[99]
  PIN state[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1239.840 2499.000 1240.400 ;
    END
  END state[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 2481.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 2481.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 2481.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 2481.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 2481.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 2481.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 2481.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 15.380 1099.040 2481.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1251.040 15.380 1252.640 2481.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1404.640 15.380 1406.240 2481.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1558.240 15.380 1559.840 2481.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1711.840 15.380 1713.440 2481.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1865.440 15.380 1867.040 2481.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2019.040 15.380 2020.640 2481.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2172.640 15.380 2174.240 2481.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2326.240 15.380 2327.840 2481.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2479.840 15.380 2481.440 2481.660 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 2481.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 2481.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 2481.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 2481.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 2481.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 2481.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 2481.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1174.240 15.380 1175.840 2481.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1327.840 15.380 1329.440 2481.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1481.440 15.380 1483.040 2481.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1635.040 15.380 1636.640 2481.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1788.640 15.380 1790.240 2481.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1942.240 15.380 1943.840 2481.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2095.840 15.380 2097.440 2481.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2249.440 15.380 2251.040 2481.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2403.040 15.380 2404.640 2481.660 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 14.710 2493.120 2483.450 ;
      LAYER Metal2 ;
        RECT 0.140 2499.300 2493.540 2499.700 ;
        RECT 0.140 2495.700 16.500 2499.300 ;
        RECT 17.660 2495.700 43.380 2499.300 ;
        RECT 44.540 2495.700 70.260 2499.300 ;
        RECT 71.420 2495.700 93.780 2499.300 ;
        RECT 94.940 2495.700 120.660 2499.300 ;
        RECT 121.820 2495.700 147.540 2499.300 ;
        RECT 148.700 2495.700 174.420 2499.300 ;
        RECT 175.580 2495.700 197.940 2499.300 ;
        RECT 199.100 2495.700 224.820 2499.300 ;
        RECT 225.980 2495.700 251.700 2499.300 ;
        RECT 252.860 2495.700 278.580 2499.300 ;
        RECT 279.740 2495.700 302.100 2499.300 ;
        RECT 303.260 2495.700 328.980 2499.300 ;
        RECT 330.140 2495.700 355.860 2499.300 ;
        RECT 357.020 2495.700 382.740 2499.300 ;
        RECT 383.900 2495.700 406.260 2499.300 ;
        RECT 407.420 2495.700 433.140 2499.300 ;
        RECT 434.300 2495.700 460.020 2499.300 ;
        RECT 461.180 2495.700 483.540 2499.300 ;
        RECT 484.700 2495.700 510.420 2499.300 ;
        RECT 511.580 2495.700 537.300 2499.300 ;
        RECT 538.460 2495.700 564.180 2499.300 ;
        RECT 565.340 2495.700 587.700 2499.300 ;
        RECT 588.860 2495.700 614.580 2499.300 ;
        RECT 615.740 2495.700 641.460 2499.300 ;
        RECT 642.620 2495.700 668.340 2499.300 ;
        RECT 669.500 2495.700 691.860 2499.300 ;
        RECT 693.020 2495.700 718.740 2499.300 ;
        RECT 719.900 2495.700 745.620 2499.300 ;
        RECT 746.780 2495.700 769.140 2499.300 ;
        RECT 770.300 2495.700 796.020 2499.300 ;
        RECT 797.180 2495.700 822.900 2499.300 ;
        RECT 824.060 2495.700 849.780 2499.300 ;
        RECT 850.940 2495.700 873.300 2499.300 ;
        RECT 874.460 2495.700 900.180 2499.300 ;
        RECT 901.340 2495.700 927.060 2499.300 ;
        RECT 928.220 2495.700 953.940 2499.300 ;
        RECT 955.100 2495.700 977.460 2499.300 ;
        RECT 978.620 2495.700 1004.340 2499.300 ;
        RECT 1005.500 2495.700 1031.220 2499.300 ;
        RECT 1032.380 2495.700 1054.740 2499.300 ;
        RECT 1055.900 2495.700 1081.620 2499.300 ;
        RECT 1082.780 2495.700 1108.500 2499.300 ;
        RECT 1109.660 2495.700 1135.380 2499.300 ;
        RECT 1136.540 2495.700 1158.900 2499.300 ;
        RECT 1160.060 2495.700 1185.780 2499.300 ;
        RECT 1186.940 2495.700 1212.660 2499.300 ;
        RECT 1213.820 2495.700 1239.540 2499.300 ;
        RECT 1240.700 2495.700 1263.060 2499.300 ;
        RECT 1264.220 2495.700 1289.940 2499.300 ;
        RECT 1291.100 2495.700 1316.820 2499.300 ;
        RECT 1317.980 2495.700 1343.700 2499.300 ;
        RECT 1344.860 2495.700 1367.220 2499.300 ;
        RECT 1368.380 2495.700 1394.100 2499.300 ;
        RECT 1395.260 2495.700 1420.980 2499.300 ;
        RECT 1422.140 2495.700 1444.500 2499.300 ;
        RECT 1445.660 2495.700 1471.380 2499.300 ;
        RECT 1472.540 2495.700 1498.260 2499.300 ;
        RECT 1499.420 2495.700 1525.140 2499.300 ;
        RECT 1526.300 2495.700 1548.660 2499.300 ;
        RECT 1549.820 2495.700 1575.540 2499.300 ;
        RECT 1576.700 2495.700 1602.420 2499.300 ;
        RECT 1603.580 2495.700 1629.300 2499.300 ;
        RECT 1630.460 2495.700 1652.820 2499.300 ;
        RECT 1653.980 2495.700 1679.700 2499.300 ;
        RECT 1680.860 2495.700 1706.580 2499.300 ;
        RECT 1707.740 2495.700 1730.100 2499.300 ;
        RECT 1731.260 2495.700 1756.980 2499.300 ;
        RECT 1758.140 2495.700 1783.860 2499.300 ;
        RECT 1785.020 2495.700 1810.740 2499.300 ;
        RECT 1811.900 2495.700 1834.260 2499.300 ;
        RECT 1835.420 2495.700 1861.140 2499.300 ;
        RECT 1862.300 2495.700 1888.020 2499.300 ;
        RECT 1889.180 2495.700 1914.900 2499.300 ;
        RECT 1916.060 2495.700 1938.420 2499.300 ;
        RECT 1939.580 2495.700 1965.300 2499.300 ;
        RECT 1966.460 2495.700 1992.180 2499.300 ;
        RECT 1993.340 2495.700 2015.700 2499.300 ;
        RECT 2016.860 2495.700 2042.580 2499.300 ;
        RECT 2043.740 2495.700 2069.460 2499.300 ;
        RECT 2070.620 2495.700 2096.340 2499.300 ;
        RECT 2097.500 2495.700 2119.860 2499.300 ;
        RECT 2121.020 2495.700 2146.740 2499.300 ;
        RECT 2147.900 2495.700 2173.620 2499.300 ;
        RECT 2174.780 2495.700 2200.500 2499.300 ;
        RECT 2201.660 2495.700 2224.020 2499.300 ;
        RECT 2225.180 2495.700 2250.900 2499.300 ;
        RECT 2252.060 2495.700 2277.780 2499.300 ;
        RECT 2278.940 2495.700 2304.660 2499.300 ;
        RECT 2305.820 2495.700 2328.180 2499.300 ;
        RECT 2329.340 2495.700 2355.060 2499.300 ;
        RECT 2356.220 2495.700 2381.940 2499.300 ;
        RECT 2383.100 2495.700 2405.460 2499.300 ;
        RECT 2406.620 2495.700 2432.340 2499.300 ;
        RECT 2433.500 2495.700 2459.220 2499.300 ;
        RECT 2460.380 2495.700 2486.100 2499.300 ;
        RECT 2487.260 2495.700 2493.540 2499.300 ;
        RECT 0.140 4.300 2493.540 2495.700 ;
        RECT 0.860 3.500 23.220 4.300 ;
        RECT 24.380 3.500 50.100 4.300 ;
        RECT 51.260 3.500 76.980 4.300 ;
        RECT 78.140 3.500 100.500 4.300 ;
        RECT 101.660 3.500 127.380 4.300 ;
        RECT 128.540 3.500 154.260 4.300 ;
        RECT 155.420 3.500 181.140 4.300 ;
        RECT 182.300 3.500 204.660 4.300 ;
        RECT 205.820 3.500 231.540 4.300 ;
        RECT 232.700 3.500 258.420 4.300 ;
        RECT 259.580 3.500 285.300 4.300 ;
        RECT 286.460 3.500 308.820 4.300 ;
        RECT 309.980 3.500 335.700 4.300 ;
        RECT 336.860 3.500 362.580 4.300 ;
        RECT 363.740 3.500 386.100 4.300 ;
        RECT 387.260 3.500 412.980 4.300 ;
        RECT 414.140 3.500 439.860 4.300 ;
        RECT 441.020 3.500 466.740 4.300 ;
        RECT 467.900 3.500 490.260 4.300 ;
        RECT 491.420 3.500 517.140 4.300 ;
        RECT 518.300 3.500 544.020 4.300 ;
        RECT 545.180 3.500 570.900 4.300 ;
        RECT 572.060 3.500 594.420 4.300 ;
        RECT 595.580 3.500 621.300 4.300 ;
        RECT 622.460 3.500 648.180 4.300 ;
        RECT 649.340 3.500 671.700 4.300 ;
        RECT 672.860 3.500 698.580 4.300 ;
        RECT 699.740 3.500 725.460 4.300 ;
        RECT 726.620 3.500 752.340 4.300 ;
        RECT 753.500 3.500 775.860 4.300 ;
        RECT 777.020 3.500 802.740 4.300 ;
        RECT 803.900 3.500 829.620 4.300 ;
        RECT 830.780 3.500 856.500 4.300 ;
        RECT 857.660 3.500 880.020 4.300 ;
        RECT 881.180 3.500 906.900 4.300 ;
        RECT 908.060 3.500 933.780 4.300 ;
        RECT 934.940 3.500 960.660 4.300 ;
        RECT 961.820 3.500 984.180 4.300 ;
        RECT 985.340 3.500 1011.060 4.300 ;
        RECT 1012.220 3.500 1037.940 4.300 ;
        RECT 1039.100 3.500 1061.460 4.300 ;
        RECT 1062.620 3.500 1088.340 4.300 ;
        RECT 1089.500 3.500 1115.220 4.300 ;
        RECT 1116.380 3.500 1142.100 4.300 ;
        RECT 1143.260 3.500 1165.620 4.300 ;
        RECT 1166.780 3.500 1192.500 4.300 ;
        RECT 1193.660 3.500 1219.380 4.300 ;
        RECT 1220.540 3.500 1246.260 4.300 ;
        RECT 1247.420 3.500 1269.780 4.300 ;
        RECT 1270.940 3.500 1296.660 4.300 ;
        RECT 1297.820 3.500 1323.540 4.300 ;
        RECT 1324.700 3.500 1347.060 4.300 ;
        RECT 1348.220 3.500 1373.940 4.300 ;
        RECT 1375.100 3.500 1400.820 4.300 ;
        RECT 1401.980 3.500 1427.700 4.300 ;
        RECT 1428.860 3.500 1451.220 4.300 ;
        RECT 1452.380 3.500 1478.100 4.300 ;
        RECT 1479.260 3.500 1504.980 4.300 ;
        RECT 1506.140 3.500 1531.860 4.300 ;
        RECT 1533.020 3.500 1555.380 4.300 ;
        RECT 1556.540 3.500 1582.260 4.300 ;
        RECT 1583.420 3.500 1609.140 4.300 ;
        RECT 1610.300 3.500 1632.660 4.300 ;
        RECT 1633.820 3.500 1659.540 4.300 ;
        RECT 1660.700 3.500 1686.420 4.300 ;
        RECT 1687.580 3.500 1713.300 4.300 ;
        RECT 1714.460 3.500 1736.820 4.300 ;
        RECT 1737.980 3.500 1763.700 4.300 ;
        RECT 1764.860 3.500 1790.580 4.300 ;
        RECT 1791.740 3.500 1817.460 4.300 ;
        RECT 1818.620 3.500 1840.980 4.300 ;
        RECT 1842.140 3.500 1867.860 4.300 ;
        RECT 1869.020 3.500 1894.740 4.300 ;
        RECT 1895.900 3.500 1921.620 4.300 ;
        RECT 1922.780 3.500 1945.140 4.300 ;
        RECT 1946.300 3.500 1972.020 4.300 ;
        RECT 1973.180 3.500 1998.900 4.300 ;
        RECT 2000.060 3.500 2022.420 4.300 ;
        RECT 2023.580 3.500 2049.300 4.300 ;
        RECT 2050.460 3.500 2076.180 4.300 ;
        RECT 2077.340 3.500 2103.060 4.300 ;
        RECT 2104.220 3.500 2126.580 4.300 ;
        RECT 2127.740 3.500 2153.460 4.300 ;
        RECT 2154.620 3.500 2180.340 4.300 ;
        RECT 2181.500 3.500 2207.220 4.300 ;
        RECT 2208.380 3.500 2230.740 4.300 ;
        RECT 2231.900 3.500 2257.620 4.300 ;
        RECT 2258.780 3.500 2284.500 4.300 ;
        RECT 2285.660 3.500 2308.020 4.300 ;
        RECT 2309.180 3.500 2334.900 4.300 ;
        RECT 2336.060 3.500 2361.780 4.300 ;
        RECT 2362.940 3.500 2388.660 4.300 ;
        RECT 2389.820 3.500 2412.180 4.300 ;
        RECT 2413.340 3.500 2439.060 4.300 ;
        RECT 2440.220 3.500 2465.940 4.300 ;
        RECT 2467.100 3.500 2492.820 4.300 ;
      LAYER Metal3 ;
        RECT 0.090 2492.820 0.700 2493.540 ;
        RECT 4.300 2492.820 2499.700 2493.540 ;
        RECT 0.090 2487.260 2499.700 2492.820 ;
        RECT 0.090 2486.100 2495.700 2487.260 ;
        RECT 2499.300 2486.100 2499.700 2487.260 ;
        RECT 0.090 2467.100 2499.700 2486.100 ;
        RECT 0.090 2465.940 0.700 2467.100 ;
        RECT 4.300 2465.940 2499.700 2467.100 ;
        RECT 0.090 2460.380 2499.700 2465.940 ;
        RECT 0.090 2459.220 2495.700 2460.380 ;
        RECT 2499.300 2459.220 2499.700 2460.380 ;
        RECT 0.090 2440.220 2499.700 2459.220 ;
        RECT 0.090 2439.060 0.700 2440.220 ;
        RECT 4.300 2439.060 2499.700 2440.220 ;
        RECT 0.090 2433.500 2499.700 2439.060 ;
        RECT 0.090 2432.340 2495.700 2433.500 ;
        RECT 2499.300 2432.340 2499.700 2433.500 ;
        RECT 0.090 2413.340 2499.700 2432.340 ;
        RECT 0.090 2412.180 0.700 2413.340 ;
        RECT 4.300 2412.180 2499.700 2413.340 ;
        RECT 0.090 2406.620 2499.700 2412.180 ;
        RECT 0.090 2405.460 2495.700 2406.620 ;
        RECT 2499.300 2405.460 2499.700 2406.620 ;
        RECT 0.090 2389.820 2499.700 2405.460 ;
        RECT 0.090 2388.660 0.700 2389.820 ;
        RECT 4.300 2388.660 2499.700 2389.820 ;
        RECT 0.090 2383.100 2499.700 2388.660 ;
        RECT 0.090 2381.940 2495.700 2383.100 ;
        RECT 2499.300 2381.940 2499.700 2383.100 ;
        RECT 0.090 2362.940 2499.700 2381.940 ;
        RECT 0.090 2361.780 0.700 2362.940 ;
        RECT 4.300 2361.780 2499.700 2362.940 ;
        RECT 0.090 2356.220 2499.700 2361.780 ;
        RECT 0.090 2355.060 2495.700 2356.220 ;
        RECT 2499.300 2355.060 2499.700 2356.220 ;
        RECT 0.090 2336.060 2499.700 2355.060 ;
        RECT 0.090 2334.900 0.700 2336.060 ;
        RECT 4.300 2334.900 2499.700 2336.060 ;
        RECT 0.090 2329.340 2499.700 2334.900 ;
        RECT 0.090 2328.180 2495.700 2329.340 ;
        RECT 2499.300 2328.180 2499.700 2329.340 ;
        RECT 0.090 2309.180 2499.700 2328.180 ;
        RECT 0.090 2308.020 0.700 2309.180 ;
        RECT 4.300 2308.020 2499.700 2309.180 ;
        RECT 0.090 2305.820 2499.700 2308.020 ;
        RECT 0.090 2304.660 2495.700 2305.820 ;
        RECT 2499.300 2304.660 2499.700 2305.820 ;
        RECT 0.090 2285.660 2499.700 2304.660 ;
        RECT 0.090 2284.500 0.700 2285.660 ;
        RECT 4.300 2284.500 2499.700 2285.660 ;
        RECT 0.090 2278.940 2499.700 2284.500 ;
        RECT 0.090 2277.780 2495.700 2278.940 ;
        RECT 2499.300 2277.780 2499.700 2278.940 ;
        RECT 0.090 2258.780 2499.700 2277.780 ;
        RECT 0.090 2257.620 0.700 2258.780 ;
        RECT 4.300 2257.620 2499.700 2258.780 ;
        RECT 0.090 2252.060 2499.700 2257.620 ;
        RECT 0.090 2250.900 2495.700 2252.060 ;
        RECT 2499.300 2250.900 2499.700 2252.060 ;
        RECT 0.090 2231.900 2499.700 2250.900 ;
        RECT 0.090 2230.740 0.700 2231.900 ;
        RECT 4.300 2230.740 2499.700 2231.900 ;
        RECT 0.090 2225.180 2499.700 2230.740 ;
        RECT 0.090 2224.020 2495.700 2225.180 ;
        RECT 2499.300 2224.020 2499.700 2225.180 ;
        RECT 0.090 2208.380 2499.700 2224.020 ;
        RECT 0.090 2207.220 0.700 2208.380 ;
        RECT 4.300 2207.220 2499.700 2208.380 ;
        RECT 0.090 2201.660 2499.700 2207.220 ;
        RECT 0.090 2200.500 2495.700 2201.660 ;
        RECT 2499.300 2200.500 2499.700 2201.660 ;
        RECT 0.090 2181.500 2499.700 2200.500 ;
        RECT 0.090 2180.340 0.700 2181.500 ;
        RECT 4.300 2180.340 2499.700 2181.500 ;
        RECT 0.090 2174.780 2499.700 2180.340 ;
        RECT 0.090 2173.620 2495.700 2174.780 ;
        RECT 2499.300 2173.620 2499.700 2174.780 ;
        RECT 0.090 2154.620 2499.700 2173.620 ;
        RECT 0.090 2153.460 0.700 2154.620 ;
        RECT 4.300 2153.460 2499.700 2154.620 ;
        RECT 0.090 2147.900 2499.700 2153.460 ;
        RECT 0.090 2146.740 2495.700 2147.900 ;
        RECT 2499.300 2146.740 2499.700 2147.900 ;
        RECT 0.090 2127.740 2499.700 2146.740 ;
        RECT 0.090 2126.580 0.700 2127.740 ;
        RECT 4.300 2126.580 2499.700 2127.740 ;
        RECT 0.090 2121.020 2499.700 2126.580 ;
        RECT 0.090 2119.860 2495.700 2121.020 ;
        RECT 2499.300 2119.860 2499.700 2121.020 ;
        RECT 0.090 2104.220 2499.700 2119.860 ;
        RECT 0.090 2103.060 0.700 2104.220 ;
        RECT 4.300 2103.060 2499.700 2104.220 ;
        RECT 0.090 2097.500 2499.700 2103.060 ;
        RECT 0.090 2096.340 2495.700 2097.500 ;
        RECT 2499.300 2096.340 2499.700 2097.500 ;
        RECT 0.090 2077.340 2499.700 2096.340 ;
        RECT 0.090 2076.180 0.700 2077.340 ;
        RECT 4.300 2076.180 2499.700 2077.340 ;
        RECT 0.090 2070.620 2499.700 2076.180 ;
        RECT 0.090 2069.460 2495.700 2070.620 ;
        RECT 2499.300 2069.460 2499.700 2070.620 ;
        RECT 0.090 2050.460 2499.700 2069.460 ;
        RECT 0.090 2049.300 0.700 2050.460 ;
        RECT 4.300 2049.300 2499.700 2050.460 ;
        RECT 0.090 2043.740 2499.700 2049.300 ;
        RECT 0.090 2042.580 2495.700 2043.740 ;
        RECT 2499.300 2042.580 2499.700 2043.740 ;
        RECT 0.090 2023.580 2499.700 2042.580 ;
        RECT 0.090 2022.420 0.700 2023.580 ;
        RECT 4.300 2022.420 2499.700 2023.580 ;
        RECT 0.090 2016.860 2499.700 2022.420 ;
        RECT 0.090 2015.700 2495.700 2016.860 ;
        RECT 2499.300 2015.700 2499.700 2016.860 ;
        RECT 0.090 2000.060 2499.700 2015.700 ;
        RECT 0.090 1998.900 0.700 2000.060 ;
        RECT 4.300 1998.900 2499.700 2000.060 ;
        RECT 0.090 1993.340 2499.700 1998.900 ;
        RECT 0.090 1992.180 2495.700 1993.340 ;
        RECT 2499.300 1992.180 2499.700 1993.340 ;
        RECT 0.090 1973.180 2499.700 1992.180 ;
        RECT 0.090 1972.020 0.700 1973.180 ;
        RECT 4.300 1972.020 2499.700 1973.180 ;
        RECT 0.090 1966.460 2499.700 1972.020 ;
        RECT 0.090 1965.300 2495.700 1966.460 ;
        RECT 2499.300 1965.300 2499.700 1966.460 ;
        RECT 0.090 1946.300 2499.700 1965.300 ;
        RECT 0.090 1945.140 0.700 1946.300 ;
        RECT 4.300 1945.140 2499.700 1946.300 ;
        RECT 0.090 1939.580 2499.700 1945.140 ;
        RECT 0.090 1938.420 2495.700 1939.580 ;
        RECT 2499.300 1938.420 2499.700 1939.580 ;
        RECT 0.090 1922.780 2499.700 1938.420 ;
        RECT 0.090 1921.620 0.700 1922.780 ;
        RECT 4.300 1921.620 2499.700 1922.780 ;
        RECT 0.090 1916.060 2499.700 1921.620 ;
        RECT 0.090 1914.900 2495.700 1916.060 ;
        RECT 2499.300 1914.900 2499.700 1916.060 ;
        RECT 0.090 1895.900 2499.700 1914.900 ;
        RECT 0.090 1894.740 0.700 1895.900 ;
        RECT 4.300 1894.740 2499.700 1895.900 ;
        RECT 0.090 1889.180 2499.700 1894.740 ;
        RECT 0.090 1888.020 2495.700 1889.180 ;
        RECT 2499.300 1888.020 2499.700 1889.180 ;
        RECT 0.090 1869.020 2499.700 1888.020 ;
        RECT 0.090 1867.860 0.700 1869.020 ;
        RECT 4.300 1867.860 2499.700 1869.020 ;
        RECT 0.090 1862.300 2499.700 1867.860 ;
        RECT 0.090 1861.140 2495.700 1862.300 ;
        RECT 2499.300 1861.140 2499.700 1862.300 ;
        RECT 0.090 1842.140 2499.700 1861.140 ;
        RECT 0.090 1840.980 0.700 1842.140 ;
        RECT 4.300 1840.980 2499.700 1842.140 ;
        RECT 0.090 1835.420 2499.700 1840.980 ;
        RECT 0.090 1834.260 2495.700 1835.420 ;
        RECT 2499.300 1834.260 2499.700 1835.420 ;
        RECT 0.090 1818.620 2499.700 1834.260 ;
        RECT 0.090 1817.460 0.700 1818.620 ;
        RECT 4.300 1817.460 2499.700 1818.620 ;
        RECT 0.090 1811.900 2499.700 1817.460 ;
        RECT 0.090 1810.740 2495.700 1811.900 ;
        RECT 2499.300 1810.740 2499.700 1811.900 ;
        RECT 0.090 1791.740 2499.700 1810.740 ;
        RECT 0.090 1790.580 0.700 1791.740 ;
        RECT 4.300 1790.580 2499.700 1791.740 ;
        RECT 0.090 1785.020 2499.700 1790.580 ;
        RECT 0.090 1783.860 2495.700 1785.020 ;
        RECT 2499.300 1783.860 2499.700 1785.020 ;
        RECT 0.090 1764.860 2499.700 1783.860 ;
        RECT 0.090 1763.700 0.700 1764.860 ;
        RECT 4.300 1763.700 2499.700 1764.860 ;
        RECT 0.090 1758.140 2499.700 1763.700 ;
        RECT 0.090 1756.980 2495.700 1758.140 ;
        RECT 2499.300 1756.980 2499.700 1758.140 ;
        RECT 0.090 1737.980 2499.700 1756.980 ;
        RECT 0.090 1736.820 0.700 1737.980 ;
        RECT 4.300 1736.820 2499.700 1737.980 ;
        RECT 0.090 1731.260 2499.700 1736.820 ;
        RECT 0.090 1730.100 2495.700 1731.260 ;
        RECT 2499.300 1730.100 2499.700 1731.260 ;
        RECT 0.090 1714.460 2499.700 1730.100 ;
        RECT 0.090 1713.300 0.700 1714.460 ;
        RECT 4.300 1713.300 2499.700 1714.460 ;
        RECT 0.090 1707.740 2499.700 1713.300 ;
        RECT 0.090 1706.580 2495.700 1707.740 ;
        RECT 2499.300 1706.580 2499.700 1707.740 ;
        RECT 0.090 1687.580 2499.700 1706.580 ;
        RECT 0.090 1686.420 0.700 1687.580 ;
        RECT 4.300 1686.420 2499.700 1687.580 ;
        RECT 0.090 1680.860 2499.700 1686.420 ;
        RECT 0.090 1679.700 2495.700 1680.860 ;
        RECT 2499.300 1679.700 2499.700 1680.860 ;
        RECT 0.090 1660.700 2499.700 1679.700 ;
        RECT 0.090 1659.540 0.700 1660.700 ;
        RECT 4.300 1659.540 2499.700 1660.700 ;
        RECT 0.090 1653.980 2499.700 1659.540 ;
        RECT 0.090 1652.820 2495.700 1653.980 ;
        RECT 2499.300 1652.820 2499.700 1653.980 ;
        RECT 0.090 1633.820 2499.700 1652.820 ;
        RECT 0.090 1632.660 0.700 1633.820 ;
        RECT 4.300 1632.660 2499.700 1633.820 ;
        RECT 0.090 1630.460 2499.700 1632.660 ;
        RECT 0.090 1629.300 2495.700 1630.460 ;
        RECT 2499.300 1629.300 2499.700 1630.460 ;
        RECT 0.090 1610.300 2499.700 1629.300 ;
        RECT 0.090 1609.140 0.700 1610.300 ;
        RECT 4.300 1609.140 2499.700 1610.300 ;
        RECT 0.090 1603.580 2499.700 1609.140 ;
        RECT 0.090 1602.420 2495.700 1603.580 ;
        RECT 2499.300 1602.420 2499.700 1603.580 ;
        RECT 0.090 1583.420 2499.700 1602.420 ;
        RECT 0.090 1582.260 0.700 1583.420 ;
        RECT 4.300 1582.260 2499.700 1583.420 ;
        RECT 0.090 1576.700 2499.700 1582.260 ;
        RECT 0.090 1575.540 2495.700 1576.700 ;
        RECT 2499.300 1575.540 2499.700 1576.700 ;
        RECT 0.090 1556.540 2499.700 1575.540 ;
        RECT 0.090 1555.380 0.700 1556.540 ;
        RECT 4.300 1555.380 2499.700 1556.540 ;
        RECT 0.090 1549.820 2499.700 1555.380 ;
        RECT 0.090 1548.660 2495.700 1549.820 ;
        RECT 2499.300 1548.660 2499.700 1549.820 ;
        RECT 0.090 1533.020 2499.700 1548.660 ;
        RECT 0.090 1531.860 0.700 1533.020 ;
        RECT 4.300 1531.860 2499.700 1533.020 ;
        RECT 0.090 1526.300 2499.700 1531.860 ;
        RECT 0.090 1525.140 2495.700 1526.300 ;
        RECT 2499.300 1525.140 2499.700 1526.300 ;
        RECT 0.090 1506.140 2499.700 1525.140 ;
        RECT 0.090 1504.980 0.700 1506.140 ;
        RECT 4.300 1504.980 2499.700 1506.140 ;
        RECT 0.090 1499.420 2499.700 1504.980 ;
        RECT 0.090 1498.260 2495.700 1499.420 ;
        RECT 2499.300 1498.260 2499.700 1499.420 ;
        RECT 0.090 1479.260 2499.700 1498.260 ;
        RECT 0.090 1478.100 0.700 1479.260 ;
        RECT 4.300 1478.100 2499.700 1479.260 ;
        RECT 0.090 1472.540 2499.700 1478.100 ;
        RECT 0.090 1471.380 2495.700 1472.540 ;
        RECT 2499.300 1471.380 2499.700 1472.540 ;
        RECT 0.090 1452.380 2499.700 1471.380 ;
        RECT 0.090 1451.220 0.700 1452.380 ;
        RECT 4.300 1451.220 2499.700 1452.380 ;
        RECT 0.090 1445.660 2499.700 1451.220 ;
        RECT 0.090 1444.500 2495.700 1445.660 ;
        RECT 2499.300 1444.500 2499.700 1445.660 ;
        RECT 0.090 1428.860 2499.700 1444.500 ;
        RECT 0.090 1427.700 0.700 1428.860 ;
        RECT 4.300 1427.700 2499.700 1428.860 ;
        RECT 0.090 1422.140 2499.700 1427.700 ;
        RECT 0.090 1420.980 2495.700 1422.140 ;
        RECT 2499.300 1420.980 2499.700 1422.140 ;
        RECT 0.090 1401.980 2499.700 1420.980 ;
        RECT 0.090 1400.820 0.700 1401.980 ;
        RECT 4.300 1400.820 2499.700 1401.980 ;
        RECT 0.090 1395.260 2499.700 1400.820 ;
        RECT 0.090 1394.100 2495.700 1395.260 ;
        RECT 2499.300 1394.100 2499.700 1395.260 ;
        RECT 0.090 1375.100 2499.700 1394.100 ;
        RECT 0.090 1373.940 0.700 1375.100 ;
        RECT 4.300 1373.940 2499.700 1375.100 ;
        RECT 0.090 1368.380 2499.700 1373.940 ;
        RECT 0.090 1367.220 2495.700 1368.380 ;
        RECT 2499.300 1367.220 2499.700 1368.380 ;
        RECT 0.090 1348.220 2499.700 1367.220 ;
        RECT 0.090 1347.060 0.700 1348.220 ;
        RECT 4.300 1347.060 2499.700 1348.220 ;
        RECT 0.090 1344.860 2499.700 1347.060 ;
        RECT 0.090 1343.700 2495.700 1344.860 ;
        RECT 2499.300 1343.700 2499.700 1344.860 ;
        RECT 0.090 1324.700 2499.700 1343.700 ;
        RECT 0.090 1323.540 0.700 1324.700 ;
        RECT 4.300 1323.540 2499.700 1324.700 ;
        RECT 0.090 1317.980 2499.700 1323.540 ;
        RECT 0.090 1316.820 2495.700 1317.980 ;
        RECT 2499.300 1316.820 2499.700 1317.980 ;
        RECT 0.090 1297.820 2499.700 1316.820 ;
        RECT 0.090 1296.660 0.700 1297.820 ;
        RECT 4.300 1296.660 2499.700 1297.820 ;
        RECT 0.090 1291.100 2499.700 1296.660 ;
        RECT 0.090 1289.940 2495.700 1291.100 ;
        RECT 2499.300 1289.940 2499.700 1291.100 ;
        RECT 0.090 1270.940 2499.700 1289.940 ;
        RECT 0.090 1269.780 0.700 1270.940 ;
        RECT 4.300 1269.780 2499.700 1270.940 ;
        RECT 0.090 1264.220 2499.700 1269.780 ;
        RECT 0.090 1263.060 2495.700 1264.220 ;
        RECT 2499.300 1263.060 2499.700 1264.220 ;
        RECT 0.090 1247.420 2499.700 1263.060 ;
        RECT 0.090 1246.260 0.700 1247.420 ;
        RECT 4.300 1246.260 2499.700 1247.420 ;
        RECT 0.090 1240.700 2499.700 1246.260 ;
        RECT 0.090 1239.540 2495.700 1240.700 ;
        RECT 2499.300 1239.540 2499.700 1240.700 ;
        RECT 0.090 1220.540 2499.700 1239.540 ;
        RECT 0.090 1219.380 0.700 1220.540 ;
        RECT 4.300 1219.380 2499.700 1220.540 ;
        RECT 0.090 1213.820 2499.700 1219.380 ;
        RECT 0.090 1212.660 2495.700 1213.820 ;
        RECT 2499.300 1212.660 2499.700 1213.820 ;
        RECT 0.090 1193.660 2499.700 1212.660 ;
        RECT 0.090 1192.500 0.700 1193.660 ;
        RECT 4.300 1192.500 2499.700 1193.660 ;
        RECT 0.090 1186.940 2499.700 1192.500 ;
        RECT 0.090 1185.780 2495.700 1186.940 ;
        RECT 2499.300 1185.780 2499.700 1186.940 ;
        RECT 0.090 1166.780 2499.700 1185.780 ;
        RECT 0.090 1165.620 0.700 1166.780 ;
        RECT 4.300 1165.620 2499.700 1166.780 ;
        RECT 0.090 1160.060 2499.700 1165.620 ;
        RECT 0.090 1158.900 2495.700 1160.060 ;
        RECT 2499.300 1158.900 2499.700 1160.060 ;
        RECT 0.090 1143.260 2499.700 1158.900 ;
        RECT 0.090 1142.100 0.700 1143.260 ;
        RECT 4.300 1142.100 2499.700 1143.260 ;
        RECT 0.090 1136.540 2499.700 1142.100 ;
        RECT 0.090 1135.380 2495.700 1136.540 ;
        RECT 2499.300 1135.380 2499.700 1136.540 ;
        RECT 0.090 1116.380 2499.700 1135.380 ;
        RECT 0.090 1115.220 0.700 1116.380 ;
        RECT 4.300 1115.220 2499.700 1116.380 ;
        RECT 0.090 1109.660 2499.700 1115.220 ;
        RECT 0.090 1108.500 2495.700 1109.660 ;
        RECT 2499.300 1108.500 2499.700 1109.660 ;
        RECT 0.090 1089.500 2499.700 1108.500 ;
        RECT 0.090 1088.340 0.700 1089.500 ;
        RECT 4.300 1088.340 2499.700 1089.500 ;
        RECT 0.090 1082.780 2499.700 1088.340 ;
        RECT 0.090 1081.620 2495.700 1082.780 ;
        RECT 2499.300 1081.620 2499.700 1082.780 ;
        RECT 0.090 1062.620 2499.700 1081.620 ;
        RECT 0.090 1061.460 0.700 1062.620 ;
        RECT 4.300 1061.460 2499.700 1062.620 ;
        RECT 0.090 1055.900 2499.700 1061.460 ;
        RECT 0.090 1054.740 2495.700 1055.900 ;
        RECT 2499.300 1054.740 2499.700 1055.900 ;
        RECT 0.090 1039.100 2499.700 1054.740 ;
        RECT 0.090 1037.940 0.700 1039.100 ;
        RECT 4.300 1037.940 2499.700 1039.100 ;
        RECT 0.090 1032.380 2499.700 1037.940 ;
        RECT 0.090 1031.220 2495.700 1032.380 ;
        RECT 2499.300 1031.220 2499.700 1032.380 ;
        RECT 0.090 1012.220 2499.700 1031.220 ;
        RECT 0.090 1011.060 0.700 1012.220 ;
        RECT 4.300 1011.060 2499.700 1012.220 ;
        RECT 0.090 1005.500 2499.700 1011.060 ;
        RECT 0.090 1004.340 2495.700 1005.500 ;
        RECT 2499.300 1004.340 2499.700 1005.500 ;
        RECT 0.090 985.340 2499.700 1004.340 ;
        RECT 0.090 984.180 0.700 985.340 ;
        RECT 4.300 984.180 2499.700 985.340 ;
        RECT 0.090 978.620 2499.700 984.180 ;
        RECT 0.090 977.460 2495.700 978.620 ;
        RECT 2499.300 977.460 2499.700 978.620 ;
        RECT 0.090 961.820 2499.700 977.460 ;
        RECT 0.090 960.660 0.700 961.820 ;
        RECT 4.300 960.660 2499.700 961.820 ;
        RECT 0.090 955.100 2499.700 960.660 ;
        RECT 0.090 953.940 2495.700 955.100 ;
        RECT 2499.300 953.940 2499.700 955.100 ;
        RECT 0.090 934.940 2499.700 953.940 ;
        RECT 0.090 933.780 0.700 934.940 ;
        RECT 4.300 933.780 2499.700 934.940 ;
        RECT 0.090 928.220 2499.700 933.780 ;
        RECT 0.090 927.060 2495.700 928.220 ;
        RECT 2499.300 927.060 2499.700 928.220 ;
        RECT 0.090 908.060 2499.700 927.060 ;
        RECT 0.090 906.900 0.700 908.060 ;
        RECT 4.300 906.900 2499.700 908.060 ;
        RECT 0.090 901.340 2499.700 906.900 ;
        RECT 0.090 900.180 2495.700 901.340 ;
        RECT 2499.300 900.180 2499.700 901.340 ;
        RECT 0.090 881.180 2499.700 900.180 ;
        RECT 0.090 880.020 0.700 881.180 ;
        RECT 4.300 880.020 2499.700 881.180 ;
        RECT 0.090 874.460 2499.700 880.020 ;
        RECT 0.090 873.300 2495.700 874.460 ;
        RECT 2499.300 873.300 2499.700 874.460 ;
        RECT 0.090 857.660 2499.700 873.300 ;
        RECT 0.090 856.500 0.700 857.660 ;
        RECT 4.300 856.500 2499.700 857.660 ;
        RECT 0.090 850.940 2499.700 856.500 ;
        RECT 0.090 849.780 2495.700 850.940 ;
        RECT 2499.300 849.780 2499.700 850.940 ;
        RECT 0.090 830.780 2499.700 849.780 ;
        RECT 0.090 829.620 0.700 830.780 ;
        RECT 4.300 829.620 2499.700 830.780 ;
        RECT 0.090 824.060 2499.700 829.620 ;
        RECT 0.090 822.900 2495.700 824.060 ;
        RECT 2499.300 822.900 2499.700 824.060 ;
        RECT 0.090 803.900 2499.700 822.900 ;
        RECT 0.090 802.740 0.700 803.900 ;
        RECT 4.300 802.740 2499.700 803.900 ;
        RECT 0.090 797.180 2499.700 802.740 ;
        RECT 0.090 796.020 2495.700 797.180 ;
        RECT 2499.300 796.020 2499.700 797.180 ;
        RECT 0.090 777.020 2499.700 796.020 ;
        RECT 0.090 775.860 0.700 777.020 ;
        RECT 4.300 775.860 2499.700 777.020 ;
        RECT 0.090 770.300 2499.700 775.860 ;
        RECT 0.090 769.140 2495.700 770.300 ;
        RECT 2499.300 769.140 2499.700 770.300 ;
        RECT 0.090 753.500 2499.700 769.140 ;
        RECT 0.090 752.340 0.700 753.500 ;
        RECT 4.300 752.340 2499.700 753.500 ;
        RECT 0.090 746.780 2499.700 752.340 ;
        RECT 0.090 745.620 2495.700 746.780 ;
        RECT 2499.300 745.620 2499.700 746.780 ;
        RECT 0.090 726.620 2499.700 745.620 ;
        RECT 0.090 725.460 0.700 726.620 ;
        RECT 4.300 725.460 2499.700 726.620 ;
        RECT 0.090 719.900 2499.700 725.460 ;
        RECT 0.090 718.740 2495.700 719.900 ;
        RECT 2499.300 718.740 2499.700 719.900 ;
        RECT 0.090 699.740 2499.700 718.740 ;
        RECT 0.090 698.580 0.700 699.740 ;
        RECT 4.300 698.580 2499.700 699.740 ;
        RECT 0.090 693.020 2499.700 698.580 ;
        RECT 0.090 691.860 2495.700 693.020 ;
        RECT 2499.300 691.860 2499.700 693.020 ;
        RECT 0.090 672.860 2499.700 691.860 ;
        RECT 0.090 671.700 0.700 672.860 ;
        RECT 4.300 671.700 2499.700 672.860 ;
        RECT 0.090 669.500 2499.700 671.700 ;
        RECT 0.090 668.340 2495.700 669.500 ;
        RECT 2499.300 668.340 2499.700 669.500 ;
        RECT 0.090 649.340 2499.700 668.340 ;
        RECT 0.090 648.180 0.700 649.340 ;
        RECT 4.300 648.180 2499.700 649.340 ;
        RECT 0.090 642.620 2499.700 648.180 ;
        RECT 0.090 641.460 2495.700 642.620 ;
        RECT 2499.300 641.460 2499.700 642.620 ;
        RECT 0.090 622.460 2499.700 641.460 ;
        RECT 0.090 621.300 0.700 622.460 ;
        RECT 4.300 621.300 2499.700 622.460 ;
        RECT 0.090 615.740 2499.700 621.300 ;
        RECT 0.090 614.580 2495.700 615.740 ;
        RECT 2499.300 614.580 2499.700 615.740 ;
        RECT 0.090 595.580 2499.700 614.580 ;
        RECT 0.090 594.420 0.700 595.580 ;
        RECT 4.300 594.420 2499.700 595.580 ;
        RECT 0.090 588.860 2499.700 594.420 ;
        RECT 0.090 587.700 2495.700 588.860 ;
        RECT 2499.300 587.700 2499.700 588.860 ;
        RECT 0.090 572.060 2499.700 587.700 ;
        RECT 0.090 570.900 0.700 572.060 ;
        RECT 4.300 570.900 2499.700 572.060 ;
        RECT 0.090 565.340 2499.700 570.900 ;
        RECT 0.090 564.180 2495.700 565.340 ;
        RECT 2499.300 564.180 2499.700 565.340 ;
        RECT 0.090 545.180 2499.700 564.180 ;
        RECT 0.090 544.020 0.700 545.180 ;
        RECT 4.300 544.020 2499.700 545.180 ;
        RECT 0.090 538.460 2499.700 544.020 ;
        RECT 0.090 537.300 2495.700 538.460 ;
        RECT 2499.300 537.300 2499.700 538.460 ;
        RECT 0.090 518.300 2499.700 537.300 ;
        RECT 0.090 517.140 0.700 518.300 ;
        RECT 4.300 517.140 2499.700 518.300 ;
        RECT 0.090 511.580 2499.700 517.140 ;
        RECT 0.090 510.420 2495.700 511.580 ;
        RECT 2499.300 510.420 2499.700 511.580 ;
        RECT 0.090 491.420 2499.700 510.420 ;
        RECT 0.090 490.260 0.700 491.420 ;
        RECT 4.300 490.260 2499.700 491.420 ;
        RECT 0.090 484.700 2499.700 490.260 ;
        RECT 0.090 483.540 2495.700 484.700 ;
        RECT 2499.300 483.540 2499.700 484.700 ;
        RECT 0.090 467.900 2499.700 483.540 ;
        RECT 0.090 466.740 0.700 467.900 ;
        RECT 4.300 466.740 2499.700 467.900 ;
        RECT 0.090 461.180 2499.700 466.740 ;
        RECT 0.090 460.020 2495.700 461.180 ;
        RECT 2499.300 460.020 2499.700 461.180 ;
        RECT 0.090 441.020 2499.700 460.020 ;
        RECT 0.090 439.860 0.700 441.020 ;
        RECT 4.300 439.860 2499.700 441.020 ;
        RECT 0.090 434.300 2499.700 439.860 ;
        RECT 0.090 433.140 2495.700 434.300 ;
        RECT 2499.300 433.140 2499.700 434.300 ;
        RECT 0.090 414.140 2499.700 433.140 ;
        RECT 0.090 412.980 0.700 414.140 ;
        RECT 4.300 412.980 2499.700 414.140 ;
        RECT 0.090 407.420 2499.700 412.980 ;
        RECT 0.090 406.260 2495.700 407.420 ;
        RECT 2499.300 406.260 2499.700 407.420 ;
        RECT 0.090 387.260 2499.700 406.260 ;
        RECT 0.090 386.100 0.700 387.260 ;
        RECT 4.300 386.100 2499.700 387.260 ;
        RECT 0.090 383.900 2499.700 386.100 ;
        RECT 0.090 382.740 2495.700 383.900 ;
        RECT 2499.300 382.740 2499.700 383.900 ;
        RECT 0.090 363.740 2499.700 382.740 ;
        RECT 0.090 362.580 0.700 363.740 ;
        RECT 4.300 362.580 2499.700 363.740 ;
        RECT 0.090 357.020 2499.700 362.580 ;
        RECT 0.090 355.860 2495.700 357.020 ;
        RECT 2499.300 355.860 2499.700 357.020 ;
        RECT 0.090 336.860 2499.700 355.860 ;
        RECT 0.090 335.700 0.700 336.860 ;
        RECT 4.300 335.700 2499.700 336.860 ;
        RECT 0.090 330.140 2499.700 335.700 ;
        RECT 0.090 328.980 2495.700 330.140 ;
        RECT 2499.300 328.980 2499.700 330.140 ;
        RECT 0.090 309.980 2499.700 328.980 ;
        RECT 0.090 308.820 0.700 309.980 ;
        RECT 4.300 308.820 2499.700 309.980 ;
        RECT 0.090 303.260 2499.700 308.820 ;
        RECT 0.090 302.100 2495.700 303.260 ;
        RECT 2499.300 302.100 2499.700 303.260 ;
        RECT 0.090 286.460 2499.700 302.100 ;
        RECT 0.090 285.300 0.700 286.460 ;
        RECT 4.300 285.300 2499.700 286.460 ;
        RECT 0.090 279.740 2499.700 285.300 ;
        RECT 0.090 278.580 2495.700 279.740 ;
        RECT 2499.300 278.580 2499.700 279.740 ;
        RECT 0.090 259.580 2499.700 278.580 ;
        RECT 0.090 258.420 0.700 259.580 ;
        RECT 4.300 258.420 2499.700 259.580 ;
        RECT 0.090 252.860 2499.700 258.420 ;
        RECT 0.090 251.700 2495.700 252.860 ;
        RECT 2499.300 251.700 2499.700 252.860 ;
        RECT 0.090 232.700 2499.700 251.700 ;
        RECT 0.090 231.540 0.700 232.700 ;
        RECT 4.300 231.540 2499.700 232.700 ;
        RECT 0.090 225.980 2499.700 231.540 ;
        RECT 0.090 224.820 2495.700 225.980 ;
        RECT 2499.300 224.820 2499.700 225.980 ;
        RECT 0.090 205.820 2499.700 224.820 ;
        RECT 0.090 204.660 0.700 205.820 ;
        RECT 4.300 204.660 2499.700 205.820 ;
        RECT 0.090 199.100 2499.700 204.660 ;
        RECT 0.090 197.940 2495.700 199.100 ;
        RECT 2499.300 197.940 2499.700 199.100 ;
        RECT 0.090 182.300 2499.700 197.940 ;
        RECT 0.090 181.140 0.700 182.300 ;
        RECT 4.300 181.140 2499.700 182.300 ;
        RECT 0.090 175.580 2499.700 181.140 ;
        RECT 0.090 174.420 2495.700 175.580 ;
        RECT 2499.300 174.420 2499.700 175.580 ;
        RECT 0.090 155.420 2499.700 174.420 ;
        RECT 0.090 154.260 0.700 155.420 ;
        RECT 4.300 154.260 2499.700 155.420 ;
        RECT 0.090 148.700 2499.700 154.260 ;
        RECT 0.090 147.540 2495.700 148.700 ;
        RECT 2499.300 147.540 2499.700 148.700 ;
        RECT 0.090 128.540 2499.700 147.540 ;
        RECT 0.090 127.380 0.700 128.540 ;
        RECT 4.300 127.380 2499.700 128.540 ;
        RECT 0.090 121.820 2499.700 127.380 ;
        RECT 0.090 120.660 2495.700 121.820 ;
        RECT 2499.300 120.660 2499.700 121.820 ;
        RECT 0.090 101.660 2499.700 120.660 ;
        RECT 0.090 100.500 0.700 101.660 ;
        RECT 4.300 100.500 2499.700 101.660 ;
        RECT 0.090 94.940 2499.700 100.500 ;
        RECT 0.090 93.780 2495.700 94.940 ;
        RECT 2499.300 93.780 2499.700 94.940 ;
        RECT 0.090 78.140 2499.700 93.780 ;
        RECT 0.090 76.980 0.700 78.140 ;
        RECT 4.300 76.980 2499.700 78.140 ;
        RECT 0.090 71.420 2499.700 76.980 ;
        RECT 0.090 70.260 2495.700 71.420 ;
        RECT 2499.300 70.260 2499.700 71.420 ;
        RECT 0.090 51.260 2499.700 70.260 ;
        RECT 0.090 50.100 0.700 51.260 ;
        RECT 4.300 50.100 2499.700 51.260 ;
        RECT 0.090 44.540 2499.700 50.100 ;
        RECT 0.090 43.380 2495.700 44.540 ;
        RECT 2499.300 43.380 2499.700 44.540 ;
        RECT 0.090 24.380 2499.700 43.380 ;
        RECT 0.090 23.220 0.700 24.380 ;
        RECT 4.300 23.220 2499.700 24.380 ;
        RECT 0.090 17.660 2499.700 23.220 ;
        RECT 0.090 16.500 2495.700 17.660 ;
        RECT 2499.300 16.500 2499.700 17.660 ;
        RECT 0.090 5.740 2499.700 16.500 ;
      LAYER Metal4 ;
        RECT 335.020 24.730 405.940 2478.470 ;
        RECT 408.140 24.730 482.740 2478.470 ;
        RECT 484.940 24.730 559.540 2478.470 ;
        RECT 561.740 24.730 636.340 2478.470 ;
        RECT 638.540 24.730 713.140 2478.470 ;
        RECT 715.340 24.730 789.940 2478.470 ;
        RECT 792.140 24.730 866.740 2478.470 ;
        RECT 868.940 24.730 943.540 2478.470 ;
        RECT 945.740 24.730 1020.340 2478.470 ;
        RECT 1022.540 24.730 1097.140 2478.470 ;
        RECT 1099.340 24.730 1173.940 2478.470 ;
        RECT 1176.140 24.730 1250.740 2478.470 ;
        RECT 1252.940 24.730 1327.540 2478.470 ;
        RECT 1329.740 24.730 1404.340 2478.470 ;
        RECT 1406.540 24.730 1481.140 2478.470 ;
        RECT 1483.340 24.730 1557.940 2478.470 ;
        RECT 1560.140 24.730 1634.740 2478.470 ;
        RECT 1636.940 24.730 1711.540 2478.470 ;
        RECT 1713.740 24.730 1788.340 2478.470 ;
        RECT 1790.540 24.730 1865.140 2478.470 ;
        RECT 1867.340 24.730 1941.940 2478.470 ;
        RECT 1944.140 24.730 2018.740 2478.470 ;
        RECT 2020.940 24.730 2095.540 2478.470 ;
        RECT 2097.740 24.730 2172.340 2478.470 ;
        RECT 2174.540 24.730 2249.140 2478.470 ;
        RECT 2251.340 24.730 2325.940 2478.470 ;
        RECT 2328.140 24.730 2402.740 2478.470 ;
        RECT 2404.940 24.730 2479.540 2478.470 ;
        RECT 2481.740 24.730 2488.500 2478.470 ;
  END
END aes128
END LIBRARY

